/* Verilog module written by vlog2Verilog (qflow) */

module mips(
    output MemRead,
    output MemWrite,
    input clk,
    output [31:0] memoryAddress,
    input [31:0] memoryOutData,
    output [31:0] memoryWriteData,
    input rst
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _6321__bF$buf0 ;
wire _6321__bF$buf1 ;
wire _6321__bF$buf2 ;
wire _6321__bF$buf3 ;
wire _6321__bF$buf4 ;
wire _5757_ ;
wire _5337_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf2  ;
wire _1677_ ;
wire [31:0] _1257_ ;
wire _7903_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _8021_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire IRWrite_bF$buf0 ;
wire _1486_ ;
wire IRWrite_bF$buf1 ;
wire _1066_ ;
wire IRWrite_bF$buf2 ;
wire IRWrite_bF$buf3 ;
wire IRWrite_bF$buf4 ;
wire _7712_ ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _8250_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _7941_ ;
wire _7521_ ;
wire _7101_ ;
wire _8306_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _7750_ ;
wire _7330_ ;
wire _8115_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _7806_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf1  ;
wire _8344_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf4  ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire [31:0] _1389_ ;
wire _7615_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _6238__bF$buf0 ;
wire _6238__bF$buf1 ;
wire _6238__bF$buf2 ;
wire _6238__bF$buf3 ;
wire _6238__bF$buf4 ;
wire _8153_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _7844_ ;
wire _7424_ ;
wire _7004_ ;
wire _8209_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _8382_ ;
wire _1830_ ;
wire _1410_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf0  ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _7653_ ;
wire _7233_ ;
wire _8018_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _8191_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf4  ;
wire _57_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf0  ;
wire _6924_ ;
wire _6504_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _7709_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _7882_ ;
wire _7462_ ;
wire _7042_ ;
wire _8247_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf4  ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf2  ;
wire _7938_ ;
wire _7518_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _7691_ ;
wire _7271_ ;
wire _8056_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf3  ;
wire _7747_ ;
wire _7327_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _7080_ ;
wire _5813_ ;
wire _8285_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf0  ;
wire _6771_ ;
wire _6351_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf3  ;
wire _7976_ ;
wire _7556_ ;
wire _7136_ ;
wire _2691_ ;
wire _2271_ ;
wire _3671__bF$buf0 ;
wire _3671__bF$buf1 ;
wire _3671__bF$buf2 ;
wire _3671__bF$buf3 ;
wire _3671__bF$buf4 ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _8094_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6580_ ;
wire _6160_ ;
wire _7785_ ;
wire _7365_ ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _7594_ ;
wire _7174_ ;
wire _5907_ ;
wire _8379_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf3  ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _8188_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _7879_ ;
wire _7459_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire [31:0] \datapath_1.regfile_1.regOut[13]  ;
wire _4177__bF$buf0 ;
wire _4177__bF$buf1 ;
wire _4177__bF$buf2 ;
wire _4177__bF$buf3 ;
wire _4177__bF$buf4 ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _7688_ ;
wire _7268_ ;
wire _3188_ ;
wire _4181__bF$buf0 ;
wire _4181__bF$buf1 ;
wire _5754_ ;
wire _4181__bF$buf2 ;
wire _5334_ ;
wire _4181__bF$buf3 ;
wire _4181__bF$buf4 ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _7900_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _7497_ ;
wire _7077_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire \datapath_1.PCJump_27_bF$buf2  ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _8303_ ;
wire _4643_ ;
wire _4223_ ;
wire [31:0] \datapath_1.regfile_1.regOut[7]  ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf2  ;
wire _8112_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _7803_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _8341_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf1  ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _7612_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _8150_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7841_ ;
wire _7421_ ;
wire _7001_ ;
wire _8206_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _7650_ ;
wire _7230_ ;
wire _8015_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf1  ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf4  ;
wire _7706_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _8244_ ;
wire _1322__bF$buf0 ;
wire _1322__bF$buf1 ;
wire _1322__bF$buf2 ;
wire _1322__bF$buf3 ;
wire _1322__bF$buf4 ;
wire _4584_ ;
wire _4164_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf1  ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _7935_ ;
wire _7515_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _8053_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf0  ;
wire _7744_ ;
wire _7324_ ;
wire _8109_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _8282_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf0  ;
wire _7973_ ;
wire _7553_ ;
wire _7133_ ;
wire _8338_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire PCWrite ;
wire _4678_ ;
wire _4258_ ;
wire _3079__bF$buf0 ;
wire _3079__bF$buf1 ;
wire _3079__bF$buf2 ;
wire _3079__bF$buf3 ;
wire _3079__bF$buf4 ;
wire _8091_ ;
wire _6824_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _7609_ ;
wire _2744_ ;
wire _2324_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf4  ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf2  ;
wire _7782_ ;
wire _7362_ ;
wire _8147_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _7838_ ;
wire _7418_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _7591_ ;
wire _7171_ ;
wire _5904_ ;
wire _8376_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire _7647_ ;
wire _7227_ ;
wire _2782_ ;
wire _2362_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf0  ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf3  ;
wire _5713_ ;
wire _8185_ ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _7876_ ;
wire _7456_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire _3796_ ;
wire _3376_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf3  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire \datapath_1.PCJump_22_bF$buf3  ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _7685_ ;
wire _7265_ ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6956_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _7494_ ;
wire _7074_ ;
wire _5807_ ;
wire _8279_ ;
wire _6264__bF$buf0 ;
wire _6264__bF$buf1 ;
wire _6264__bF$buf2 ;
wire _6264__bF$buf3 ;
wire _6264__bF$buf4 ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf3  ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _8088_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire _7779_ ;
wire _7359_ ;
wire _2494_ ;
wire _2074_ ;
wire _8300_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _7588_ ;
wire _7168_ ;
wire _3737__bF$buf0 ;
wire _3737__bF$buf1 ;
wire _3737__bF$buf2 ;
wire _3737__bF$buf3 ;
wire _3737__bF$buf4 ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _7800_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _7397_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf2  ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire _8203_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf2  ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _8012_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf1  ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _7703_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _8241_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _7932_ ;
wire _7512_ ;
wire _197_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _8050_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _7741_ ;
wire _7321_ ;
wire _8106_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf1  ;
wire _3717_ ;
wire _6189_ ;
wire _7970_ ;
wire _7550_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf4  ;
wire _7130_ ;
wire _8335_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _7606_ ;
wire _2741_ ;
wire _2321_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf1  ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf4  ;
wire _7_ ;
wire _8144_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _7835_ ;
wire _7415_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _8373_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _1916__bF$buf0 ;
wire _1916__bF$buf1 ;
wire _1916__bF$buf2 ;
wire _732_ ;
wire _1916__bF$buf3 ;
wire _312_ ;
wire _1916__bF$buf4 ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _7644_ ;
wire _7224_ ;
wire _2048__bF$buf0 ;
wire _2048__bF$buf1 ;
wire _2048__bF$buf2 ;
wire _2048__bF$buf3 ;
wire _2048__bF$buf4 ;
wire _8009_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf0  ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _8182_ ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _7873_ ;
wire _7453_ ;
wire _7033_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf4  ;
wire _8238_ ;
wire _3793_ ;
wire _3373_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf0  ;
wire _4998_ ;
wire _4578_ ;
wire Branch ;
wire _4158_ ;
wire \datapath_1.PCJump_22_bF$buf0  ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _7929_ ;
wire _7509_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _7682_ ;
wire _7262_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf4  ;
wire _8047_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire _7738_ ;
wire _7318_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _7491_ ;
wire _7071_ ;
wire _5804_ ;
wire _8276_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf3  ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf0  ;
wire _6762_ ;
wire _6342_ ;
wire _7967_ ;
wire _7547_ ;
wire _7127_ ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf4  ;
wire _5613_ ;
wire _8085_ ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire _7776_ ;
wire _7356_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6315__bF$buf0 ;
wire _6315__bF$buf1 ;
wire _6315__bF$buf2 ;
wire _6315__bF$buf3 ;
wire _6315__bF$buf4 ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire rst_bF$buf110 ;
wire rst_bF$buf111 ;
wire rst_bF$buf112 ;
wire rst_bF$buf113 ;
wire _7585_ ;
wire _7165_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire [31:0] _729_ ;
wire _309_ ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _7394_ ;
wire _5707_ ;
wire _8179_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6271__bF$buf0 ;
wire _6271__bF$buf1 ;
wire _6271__bF$buf2 ;
wire _6271__bF$buf3 ;
wire _6271__bF$buf4 ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire RegDst ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _7679_ ;
wire _7259_ ;
wire _2394_ ;
wire _8200_ ;
wire _4187__bF$buf0 ;
wire _4187__bF$buf1 ;
wire _4187__bF$buf2 ;
wire _4187__bF$buf3 ;
wire _4187__bF$buf4 ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _7488_ ;
wire _7068_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _7700_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire clk_bF$buf80 ;
wire clk_bF$buf81 ;
wire clk_bF$buf82 ;
wire clk_bF$buf83 ;
wire clk_bF$buf84 ;
wire clk_bF$buf85 ;
wire _3620_ ;
wire clk_bF$buf86 ;
wire _3200_ ;
wire clk_bF$buf87 ;
wire clk_bF$buf88 ;
wire clk_bF$buf89 ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _7297_ ;
wire _5783_ ;
wire _5363_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf2  ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _8103_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf1  ;
wire _4919_ ;
wire _8332_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _7603_ ;
wire _288_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf1  ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _8141_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _7832_ ;
wire _7412_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _8370_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _7641_ ;
wire _7221_ ;
wire _8006_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _6912_ ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire _7870_ ;
wire _7450_ ;
wire _7030_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf1  ;
wire _8235_ ;
wire _3790_ ;
wire _3370_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf4  ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _7926_ ;
wire _7506_ ;
wire _2641_ ;
wire _2221_ ;
wire _4135__bF$buf0 ;
wire _4135__bF$buf1 ;
wire _4135__bF$buf2 ;
wire _4135__bF$buf3 ;
wire _4135__bF$buf4 ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf1  ;
wire _8044_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _7735_ ;
wire _7315_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _1190__bF$buf0 ;
wire _1190__bF$buf1 ;
wire _1190__bF$buf2 ;
wire _1190__bF$buf3 ;
wire _1190__bF$buf4 ;
wire _3655_ ;
wire _3235_ ;
wire _6255__bF$buf0 ;
wire _6255__bF$buf1 ;
wire _6255__bF$buf2 ;
wire _6255__bF$buf3 ;
wire _6255__bF$buf4 ;
wire _5801_ ;
wire _8273_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf0  ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _7964_ ;
wire _7544_ ;
wire _7124_ ;
wire _8329_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf1  ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _8082_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf4  ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire [31:0] _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _7773_ ;
wire _7353_ ;
wire _3089__bF$buf0 ;
wire _3089__bF$buf1 ;
wire _3089__bF$buf2 ;
wire _3089__bF$buf3 ;
wire _3089__bF$buf4 ;
wire _8138_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _7829_ ;
wire _7409_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _7582_ ;
wire _7162_ ;
wire _8367_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire _7638_ ;
wire _7218_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _7391_ ;
wire _5704_ ;
wire _8176_ ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _7867_ ;
wire _7447_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire _7676_ ;
wire _7256_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire [31:0] _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf2  ;
wire _7485_ ;
wire _7065_ ;
wire [31:0] \datapath_1.regfile_1.regOut[2]  ;
wire _662__bF$buf0 ;
wire _662__bF$buf1 ;
wire _662__bF$buf2 ;
wire _662__bF$buf3 ;
wire _662__bF$buf4 ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _7294_ ;
wire _5607_ ;
wire _8079_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf2  ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _7999_ ;
wire _7579_ ;
wire _7159_ ;
wire _2294_ ;
wire _8100_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire [31:0] \datapath_1.regfile_1.regOut[25]  ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire _7388_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _7600_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf2  ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire [31:0] _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _7197_ ;
wire _1982__bF$buf0 ;
wire _1982__bF$buf1 ;
wire _1982__bF$buf2 ;
wire _1982__bF$buf3 ;
wire _1982__bF$buf4 ;
wire _5683_ ;
wire _5263_ ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf2  ;
wire _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _8003_ ;
wire _4763_ ;
wire _4343_ ;
wire rst_bF$buf0 ;
wire rst_bF$buf1 ;
wire rst_bF$buf2 ;
wire rst_bF$buf3 ;
wire rst_bF$buf4 ;
wire _5968_ ;
wire rst_bF$buf5 ;
wire _5548_ ;
wire rst_bF$buf6 ;
wire _5128_ ;
wire rst_bF$buf7 ;
wire rst_bF$buf8 ;
wire rst_bF$buf9 ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _8232_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf1  ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _7923_ ;
wire _7503_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf2  ;
wire _4628_ ;
wire _4208_ ;
wire _8041_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _7732_ ;
wire _7312_ ;
wire _3652_ ;
wire _3232_ ;
wire _464__bF$buf0 ;
wire _464__bF$buf1 ;
wire _464__bF$buf2 ;
wire _464__bF$buf3 ;
wire _464__bF$buf4 ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _8270_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _7961_ ;
wire _7541_ ;
wire _7121_ ;
wire _8326_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf1  ;
wire _6812_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf4  ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _7770_ ;
wire _7350_ ;
wire _8135_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf4  ;
wire _7826_ ;
wire _7406_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _8364_ ;
wire _4142__bF$buf0 ;
wire _4142__bF$buf1 ;
wire _4142__bF$buf2 ;
wire _4142__bF$buf3 ;
wire _4142__bF$buf4 ;
wire _1812_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire _7635_ ;
wire _7215_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire rst_bF$buf90 ;
wire rst_bF$buf91 ;
wire rst_bF$buf92 ;
wire rst_bF$buf93 ;
wire rst_bF$buf94 ;
wire rst_bF$buf95 ;
wire rst_bF$buf96 ;
wire rst_bF$buf97 ;
wire rst_bF$buf98 ;
wire rst_bF$buf99 ;
wire _5701_ ;
wire _8173_ ;
wire _39_ ;
wire _6906_ ;
wire _6262__bF$buf0 ;
wire _6262__bF$buf1 ;
wire _6262__bF$buf2 ;
wire _6262__bF$buf3 ;
wire _6262__bF$buf4 ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _7864_ ;
wire _7444_ ;
wire _7024_ ;
wire _8229_ ;
wire _3784_ ;
wire _3364_ ;
wire _1784__bF$buf0 ;
wire _1784__bF$buf1 ;
wire _1784__bF$buf2 ;
wire _1784__bF$buf3 ;
wire _1784__bF$buf4 ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire IorD ;
wire _7673_ ;
wire _7253_ ;
wire clk ;
wire _8038_ ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _7729_ ;
wire _7309_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _7482_ ;
wire _7062_ ;
wire _8267_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _7958_ ;
wire _7538_ ;
wire _7118_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _7291_ ;
wire _5604_ ;
wire _8076_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire _7767_ ;
wire _1256__bF$buf0 ;
wire _7347_ ;
wire _1256__bF$buf1 ;
wire _1256__bF$buf2 ;
wire _1256__bF$buf3 ;
wire _1256__bF$buf4 ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _7996_ ;
wire _7576_ ;
wire _7156_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf2  ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _7385_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _7194_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _6206__bF$buf0 ;
wire _6206__bF$buf1 ;
wire _6206__bF$buf2 ;
wire _6206__bF$buf3 ;
wire _6206__bF$buf4 ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _4197__bF$buf0 ;
wire _4197__bF$buf1 ;
wire _4197__bF$buf2 ;
wire _4197__bF$buf3 ;
wire _4197__bF$buf4 ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _7899_ ;
wire _7479_ ;
wire _7059_ ;
wire _2194_ ;
wire _8000_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire [31:0] \datapath_1.regfile_1.regOut[15]  ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf4  ;
wire _4816_ ;
wire _7288_ ;
wire _5774_ ;
wire _5354_ ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _7920_ ;
wire _7500_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire _7097_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf2  ;
wire _5583_ ;
wire _5163_ ;
wire _4130__bF$buf0 ;
wire _4130__bF$buf1 ;
wire _4130__bF$buf2 ;
wire _4130__bF$buf3 ;
wire _4130__bF$buf4 ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _8323_ ;
wire _4663_ ;
wire _4243_ ;
wire [31:0] \datapath_1.regfile_1.regOut[9]  ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf1  ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _8132_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf2  ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf1  ;
wire _1597_ ;
wire _1177_ ;
wire _7823_ ;
wire _7403_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _8361_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _7632_ ;
wire _7212_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire rst_bF$buf60 ;
wire rst_bF$buf61 ;
wire rst_bF$buf62 ;
wire rst_bF$buf63 ;
wire rst_bF$buf64 ;
wire rst_bF$buf65 ;
wire rst_bF$buf66 ;
wire rst_bF$buf67 ;
wire rst_bF$buf68 ;
wire rst_bF$buf69 ;
wire _4757_ ;
wire _4337_ ;
wire _8170_ ;
wire _36_ ;
wire _6903_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _7861_ ;
wire _7441_ ;
wire _7021_ ;
wire _8226_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire _7917_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _7670_ ;
wire _7250_ ;
wire _8035_ ;
wire RegWrite ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _7726_ ;
wire _7306_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _2376__bF$buf0 ;
wire _2376__bF$buf1 ;
wire _2376__bF$buf2 ;
wire _2376__bF$buf3 ;
wire _8264_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _7955_ ;
wire _7535_ ;
wire _7115_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf3  ;
wire _5601_ ;
wire _8073_ ;
wire [31:0] \datapath_1.mux_pcsrc.dout  ;
wire _6806_ ;
wire _1941_ ;
wire [31:0] _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _7764_ ;
wire _7344_ ;
wire _8129_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _7993_ ;
wire _7573_ ;
wire _7153_ ;
wire _8358_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _7629_ ;
wire _7209_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _7382_ ;
wire _8167_ ;
wire [31:0] \datapath_1.regfile_1.regOut[30]  ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _7858_ ;
wire _7438_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire [5:0] \control_1.op  ;
wire _3778_ ;
wire _3358_ ;
wire _7191_ ;
wire _4208__bF$buf0 ;
wire _4208__bF$buf1 ;
wire _4208__bF$buf2 ;
wire _4208__bF$buf3 ;
wire _4208__bF$buf4 ;
wire _5924_ ;
wire _5504_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf2  ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire _7667_ ;
wire _7247_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6328__bF$buf0 ;
wire _6328__bF$buf1 ;
wire _6328__bF$buf2 ;
wire _6328__bF$buf3 ;
wire _6328__bF$buf4 ;
wire _6938_ ;
wire _6518_ ;
wire [31:0] _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7896_ ;
wire _7476_ ;
wire _7056_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf1  ;
wire _4813_ ;
wire _7285_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _4622_ ;
wire _4202_ ;
wire _7094_ ;
wire _5827_ ;
wire _5407_ ;
wire _8299_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf2  ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf3  ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _7799_ ;
wire _7379_ ;
wire _2094_ ;
wire [31:0] _8320_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf4  ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire [31:0] _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _7188_ ;
wire _5674_ ;
wire _5254_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf2  ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _7820_ ;
wire _7400_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf2  ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire rst_bF$buf30 ;
wire rst_bF$buf31 ;
wire rst_bF$buf32 ;
wire rst_bF$buf33 ;
wire rst_bF$buf34 ;
wire rst_bF$buf35 ;
wire rst_bF$buf36 ;
wire rst_bF$buf37 ;
wire rst_bF$buf38 ;
wire rst_bF$buf39 ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _6900_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _8223_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire _7914_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf2  ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _8032_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _7723_ ;
wire _7303_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _8261_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _7952_ ;
wire _7532_ ;
wire _7112_ ;
wire _8317_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf0  ;
wire _4657_ ;
wire _4237_ ;
wire _8070_ ;
wire _6803_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _7761_ ;
wire _7341_ ;
wire _8126_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _7817_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire _7990_ ;
wire _7570_ ;
wire _7150_ ;
wire _8355_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _2379__bF$buf0 ;
wire _2379__bF$buf1 ;
wire _2379__bF$buf2 ;
wire _2379__bF$buf3 ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire _7626_ ;
wire _7206_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _8164_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf3  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7855_ ;
wire _7435_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _6272__bF$buf0 ;
wire _6272__bF$buf1 ;
wire _6272__bF$buf2 ;
wire _6272__bF$buf3 ;
wire _6272__bF$buf4 ;
wire _5921_ ;
wire _5501_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf2  ;
wire _7664_ ;
wire _7244_ ;
wire _8029_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire [31:0] \datapath_1.Data  ;
wire _7893_ ;
wire _7473_ ;
wire _7053_ ;
wire _8258_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _7949_ ;
wire _7529_ ;
wire _7109_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _7282_ ;
wire _3350__bF$buf0 ;
wire _3350__bF$buf1 ;
wire _3350__bF$buf2 ;
wire _3350__bF$buf3 ;
wire _3350__bF$buf4 ;
wire _8067_ ;
wire [31:0] \datapath_1.regfile_1.regOut[20]  ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _7758_ ;
wire _7338_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf2  ;
wire _3678_ ;
wire _3258_ ;
wire _7091_ ;
wire _5824_ ;
wire _5404_ ;
wire _8296_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _7987_ ;
wire _7567_ ;
wire _7147_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf0  ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _7796_ ;
wire _7376_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf1  ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _6287__bF$buf0 ;
wire _6287__bF$buf1 ;
wire _6287__bF$buf2 ;
wire _6287__bF$buf3 ;
wire _6287__bF$buf4 ;
wire _4713_ ;
wire _7185_ ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf2  ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _8199_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf3  ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _6216__bF$buf0 ;
wire _6216__bF$buf1 ;
wire _6216__bF$buf2 ;
wire _6216__bF$buf3 ;
wire _6216__bF$buf4 ;
wire _2185_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire MemRead ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _7699_ ;
wire _7279_ ;
wire _8220_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _7911_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire \datapath_1.PCJump_17_bF$buf4  ;
wire _4616_ ;
wire _7088_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _7720_ ;
wire _7300_ ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _4234__bF$buf0 ;
wire _4234__bF$buf1 ;
wire _4234__bF$buf2 ;
wire _4234__bF$buf3 ;
wire _4234__bF$buf4 ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire clk_hier0_bF$buf8 ;
wire clk_hier0_bF$buf9 ;
wire _2088_ ;
wire _8314_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire _8123_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf4  ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire _7814_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _8352_ ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _7623_ ;
wire _7203_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _8161_ ;
wire _27_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf0  ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire clk_bF$buf110 ;
wire clk_bF$buf111 ;
wire clk_bF$buf112 ;
wire clk_bF$buf113 ;
wire _7852_ ;
wire _7432_ ;
wire _7012_ ;
wire _8217_ ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _6703_ ;
wire _7908_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _7661_ ;
wire _7241_ ;
wire _8026_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _7717_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf3  ;
wire _3637_ ;
wire _3217_ ;
wire _7890_ ;
wire _7470_ ;
wire _7050_ ;
wire _8255_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf3  ;
wire _7946_ ;
wire _7526_ ;
wire _7106_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _8064_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _7755_ ;
wire _7335_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf2  ;
wire _5821_ ;
wire _5401_ ;
wire _8293_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _7984_ ;
wire _7564_ ;
wire _7144_ ;
wire _8349_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _398__bF$buf0 ;
wire _398__bF$buf1 ;
wire _398__bF$buf2 ;
wire _398__bF$buf3 ;
wire _2755_ ;
wire _398__bF$buf4 ;
wire _2335_ ;
wire _4901_ ;
wire _7793_ ;
wire _7373_ ;
wire _8158_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _690_ ;
wire _270_ ;
wire _7849_ ;
wire _7429_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _7182_ ;
wire _5915_ ;
wire _8387_ ;
wire [31:0] \datapath_1.regfile_1.regOut[10]  ;
wire \datapath_1.regfile_1.regEn_18_bF$buf2  ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire _7658_ ;
wire _7238_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf2  ;
wire _5724_ ;
wire _5304_ ;
wire _8196_ ;
wire _6929_ ;
wire _6509_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf0  ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire [31:0] _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _7887_ ;
wire _7467_ ;
wire _7047_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _7696_ ;
wire _7276_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire \datapath_1.PCJump_17_bF$buf1  ;
wire _4613_ ;
wire _7085_ ;
wire [31:0] \datapath_1.regfile_1.regOut[4]  ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf3  ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _8099_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _8311_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire [31:0] _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _4707_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf4  ;
wire _7599_ ;
wire _7179_ ;
wire _8120_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf1  ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire [31:0] \datapath_1.regfile_1.regOut[27]  ;
wire _1585_ ;
wire _1165_ ;
wire _7811_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _7620_ ;
wire _7200_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire _4241__bF$buf0 ;
wire _4241__bF$buf1 ;
wire _4241__bF$buf2 ;
wire _4241__bF$buf3 ;
wire _4241__bF$buf4 ;
wire _8214_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf4  ;
wire _1679_ ;
wire _1259_ ;
wire _7905_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _8023_ ;
wire _2157__bF$buf0 ;
wire _2157__bF$buf1 ;
wire _2157__bF$buf2 ;
wire _2157__bF$buf3 ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _7714_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf0  ;
wire [31:0] _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _8252_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf0  ;
wire _1297_ ;
wire _7943_ ;
wire _7523_ ;
wire _7103_ ;
wire _8308_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _8061_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _7752_ ;
wire _7332_ ;
wire _8117_ ;
wire [31:0] _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _8290_ ;
wire _6603_ ;
wire _7808_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _7981_ ;
wire _7561_ ;
wire _7141_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf3  ;
wire _8346_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _4158__bF$buf0 ;
wire _4158__bF$buf1 ;
wire _4158__bF$buf2 ;
wire _4158__bF$buf3 ;
wire _6832_ ;
wire _4158__bF$buf4 ;
wire _6412_ ;
wire _7617_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _7790_ ;
wire _7370_ ;
wire _8155_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire MemToReg ;
wire _6641_ ;
wire _6221_ ;
wire _7846_ ;
wire _7426_ ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _8384_ ;
wire _1832_ ;
wire _1412_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf2  ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire _6282__bF$buf0 ;
wire _6282__bF$buf1 ;
wire _6282__bF$buf2 ;
wire _6282__bF$buf3 ;
wire _6282__bF$buf4 ;
wire _7655_ ;
wire _7235_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _200__bF$buf0 ;
wire _200__bF$buf1 ;
wire _200__bF$buf2 ;
wire _200__bF$buf3 ;
wire _200__bF$buf4 ;
wire _5721_ ;
wire _5301_ ;
wire _8193_ ;
wire _59_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf2  ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _7884_ ;
wire _7464_ ;
wire _7044_ ;
wire _8249_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf4  ;
wire _6211__bF$buf0 ;
wire _6211__bF$buf1 ;
wire _6211__bF$buf2 ;
wire _6211__bF$buf3 ;
wire _6211__bF$buf4 ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _7693_ ;
wire _7273_ ;
wire _8058_ ;
wire _3193_ ;
wire [31:0] \datapath_1.rd1  ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _7749_ ;
wire _7329_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _7082_ ;
wire _5815_ ;
wire _8287_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf2  ;
wire _6773_ ;
wire _6353_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf0  ;
wire _7978_ ;
wire _7558_ ;
wire _7138_ ;
wire _2693_ ;
wire _2273_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _4225__bF$buf0 ;
wire _4225__bF$buf1 ;
wire _4225__bF$buf2 ;
wire _4225__bF$buf3 ;
wire _4225__bF$buf4 ;
wire _5624_ ;
wire _5204_ ;
wire _8096_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire [5:0] \aluControl_1.inst  ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _7787_ ;
wire _7367_ ;
wire _2082_ ;
wire _3287_ ;
wire _1520__bF$buf0 ;
wire _1520__bF$buf1 ;
wire _1520__bF$buf2 ;
wire _1520__bF$buf3 ;
wire _5853_ ;
wire _1520__bF$buf4 ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf1  ;
wire _7596_ ;
wire _7176_ ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6297__bF$buf0 ;
wire _6297__bF$buf1 ;
wire _6297__bF$buf2 ;
wire _6867_ ;
wire _6297__bF$buf3 ;
wire _6447_ ;
wire _6297__bF$buf4 ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire PCEn_bF$buf0 ;
wire PCEn_bF$buf1 ;
wire PCEn_bF$buf2 ;
wire PCEn_bF$buf3 ;
wire PCEn_bF$buf4 ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _8211_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf1  ;
wire _1676_ ;
wire _1256_ ;
wire _7902_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _7499_ ;
wire _7079_ ;
wire _8020_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire [31:0] \datapath_1.regfile_1.regOut[17]  ;
wire _1485_ ;
wire _1065_ ;
wire _7711_ ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4146__bF$buf0 ;
wire _4146__bF$buf1 ;
wire _4146__bF$buf2 ;
wire _4146__bF$buf3 ;
wire _4146__bF$buf4 ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _7940_ ;
wire _7520_ ;
wire _7100_ ;
wire _2499_ ;
wire _2079_ ;
wire _8305_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf4  ;
wire _8114_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _7805_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf0  ;
wire _8343_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf3  ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _7614_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _8152_ ;
wire _3344__bF$buf0 ;
wire _3344__bF$buf1 ;
wire _3344__bF$buf2 ;
wire _3344__bF$buf3 ;
wire _3344__bF$buf4 ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7843_ ;
wire _7423_ ;
wire _7003_ ;
wire _8208_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _8381_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _7652_ ;
wire _7232_ ;
wire _8017_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _3935__bF$buf0 ;
wire _3935__bF$buf1 ;
wire _3935__bF$buf2 ;
wire _4777_ ;
wire _3935__bF$buf3 ;
wire _4357_ ;
wire _3935__bF$buf4 ;
wire _8190_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf3  ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire _7708_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _7881_ ;
wire _7461_ ;
wire _7041_ ;
wire _8246_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf3  ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf1  ;
wire _7937_ ;
wire _7517_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _7690_ ;
wire _7270_ ;
wire _8055_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf2  ;
wire _7746_ ;
wire _7326_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire [31:0] \datapath_1.alu_1.ALUInB  ;
wire _8284_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf2  ;
wire _7975_ ;
wire _7555_ ;
wire _7135_ ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _8093_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf4  ;
wire _7784_ ;
wire _7364_ ;
wire _8149_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire [3:0] \control_1.reg_state.dout  ;
wire _4701_ ;
wire _7593_ ;
wire _7173_ ;
wire _6312__bF$buf0 ;
wire _6312__bF$buf1 ;
wire _6312__bF$buf2 ;
wire _6312__bF$buf3 ;
wire _6312__bF$buf4 ;
wire _5906_ ;
wire _8378_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire _7649_ ;
wire _7229_ ;
wire _2784_ ;
wire _2364_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf2  ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _8187_ ;
wire _1635_ ;
wire _1215_ ;
wire _4228__bF$buf0 ;
wire _4228__bF$buf1 ;
wire _4228__bF$buf2 ;
wire _4228__bF$buf3 ;
wire _4228__bF$buf4 ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _7878_ ;
wire _7458_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _7687_ ;
wire _7267_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6958_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _7496_ ;
wire _7076_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire \datapath_1.PCJump_27_bF$buf1  ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _6229__bF$buf0 ;
wire _6229__bF$buf1 ;
wire _6229__bF$buf2 ;
wire _6229__bF$buf3 ;
wire _6229__bF$buf4 ;
wire _2496_ ;
wire _2076_ ;
wire _8302_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf1  ;
wire _8111_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _7802_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire _7399_ ;
wire _8340_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf0  ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _7611_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf4  ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7840_ ;
wire _7420_ ;
wire _7000_ ;
wire _2399_ ;
wire _8205_ ;
wire _3760_ ;
wire _3340_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf4  ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _8014_ ;
wire _4774_ ;
wire _4354_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf0  ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf3  ;
wire _1899_ ;
wire _1479_ ;
wire [31:0] _1059_ ;
wire _7705_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _8243_ ;
wire _4583_ ;
wire _4163_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf0  ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire _3347__bF$buf0 ;
wire _3347__bF$buf1 ;
wire _3347__bF$buf2 ;
wire _3347__bF$buf3 ;
wire _3347__bF$buf4 ;
wire _1288_ ;
wire _7934_ ;
wire _7514_ ;
wire _199_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _8052_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _6300__bF$buf0 ;
wire _6300__bF$buf1 ;
wire _6300__bF$buf2 ;
wire _5597_ ;
wire _6300__bF$buf3 ;
wire _5177_ ;
wire _6300__bF$buf4 ;
wire _91_ ;
wire _1097_ ;
wire _7743_ ;
wire _7323_ ;
wire _8108_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _8281_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf3  ;
wire _3719_ ;
wire _7972_ ;
wire _7552_ ;
wire _7132_ ;
wire _8337_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _8090_ ;
wire _6823_ ;
wire _6403_ ;
wire _7608_ ;
wire _2743_ ;
wire _2323_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf3  ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf1  ;
wire _7781_ ;
wire _7361_ ;
wire _8146_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _7837_ ;
wire _7417_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _7590_ ;
wire _7170_ ;
wire _5903_ ;
wire _4172__bF$buf0 ;
wire _4172__bF$buf1 ;
wire _4172__bF$buf2 ;
wire _4172__bF$buf3 ;
wire _4172__bF$buf4 ;
wire _8375_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire _7646_ ;
wire _7226_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf2  ;
wire _5712_ ;
wire _8184_ ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7875_ ;
wire _7455_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf2  ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire \datapath_1.PCJump_22_bF$buf2  ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _7684_ ;
wire _7264_ ;
wire _8049_ ;
wire _3184_ ;
wire _6221__bF$buf0 ;
wire _6221__bF$buf1 ;
wire _6221__bF$buf2 ;
wire [31:0] _1917_ ;
wire _6221__bF$buf3 ;
wire _6221__bF$buf4 ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6955_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _7493_ ;
wire _7073_ ;
wire _5806_ ;
wire _8278_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf2  ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _7969_ ;
wire _7549_ ;
wire _7129_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _8087_ ;
wire [31:0] \datapath_1.regfile_1.regOut[22]  ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _7778_ ;
wire _7358_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _7587_ ;
wire _7167_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _7396_ ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf1  ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire [31:0] _1191_ ;
wire _2396_ ;
wire _8202_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf1  ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _6236__bF$buf0 ;
wire _6236__bF$buf1 ;
wire _6236__bF$buf2 ;
wire _6236__bF$buf3 ;
wire _6236__bF$buf4 ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _8011_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf0  ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _7702_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _7299_ ;
wire _8240_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf4  ;
wire _1285_ ;
wire _7931_ ;
wire _7511_ ;
wire _196_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2387__bF$buf0 ;
wire _2387__bF$buf1 ;
wire _2387__bF$buf2 ;
wire _2387__bF$buf3 ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _7740_ ;
wire _7320_ ;
wire _2299_ ;
wire _8105_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf0  ;
wire _3716_ ;
wire _6188_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf3  ;
wire _8334_ ;
wire _4674_ ;
wire _4254_ ;
wire _860__bF$buf0 ;
wire _860__bF$buf1 ;
wire _860__bF$buf2 ;
wire _860__bF$buf3 ;
wire _860__bF$buf4 ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _7605_ ;
wire _2740_ ;
wire _2320_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf0  ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf3  ;
wire _6_ ;
wire _8143_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire _7834_ ;
wire _7414_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _8372_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire _7643_ ;
wire _7223_ ;
wire _8008_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _8181_ ;
wire _47_ ;
wire _6914_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire _7872_ ;
wire _7452_ ;
wire _7032_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf3  ;
wire _8237_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _7928_ ;
wire _7508_ ;
wire _2643_ ;
wire _2223_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _7681_ ;
wire _7261_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf3  ;
wire _8046_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _4175__bF$buf0 ;
wire _4175__bF$buf1 ;
wire _4175__bF$buf2 ;
wire _4175__bF$buf3 ;
wire _4175__bF$buf4 ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _7737_ ;
wire _7317_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _7490_ ;
wire _7070_ ;
wire _5803_ ;
wire _8275_ ;
wire _1723_ ;
wire _1303_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf2  ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _7966_ ;
wire _7546_ ;
wire _7126_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf3  ;
wire _5612_ ;
wire _8084_ ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire _7775_ ;
wire _7355_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire rst_bF$buf100 ;
wire rst_bF$buf101 ;
wire rst_bF$buf102 ;
wire rst_bF$buf103 ;
wire rst_bF$buf104 ;
wire rst_bF$buf105 ;
wire rst_bF$buf106 ;
wire rst_bF$buf107 ;
wire rst_bF$buf108 ;
wire rst_bF$buf109 ;
wire _7584_ ;
wire _7164_ ;
wire _8369_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _4921_ ;
wire _4501_ ;
wire _7393_ ;
wire _5706_ ;
wire _8178_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire rst ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _7869_ ;
wire _7449_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire [31:0] \datapath_1.regfile_1.regOut[12]  ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _7678_ ;
wire _7258_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf4  ;
wire MemWrite ;
wire _7487_ ;
wire _7067_ ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire clk_bF$buf76 ;
wire _134__bF$buf0 ;
wire clk_bF$buf77 ;
wire _134__bF$buf1 ;
wire clk_bF$buf78 ;
wire _134__bF$buf2 ;
wire clk_bF$buf79 ;
wire _134__bF$buf3 ;
wire _134__bF$buf4 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _7296_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf1  ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf4  ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire [31:0] \datapath_1.regfile_1.regOut[6]  ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _8102_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf0  ;
wire _4918_ ;
wire _8331_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _7602_ ;
wire _287_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf4  ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf0  ;
wire [31:0] _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _7199_ ;
wire _8140_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [31:0] \datapath_1.regfile_1.regOut[29]  ;
wire _1185_ ;
wire _7831_ ;
wire _7411_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf4  ;
wire _3751_ ;
wire _3331_ ;
wire _1454__bF$buf0 ;
wire _1454__bF$buf1 ;
wire _1454__bF$buf2 ;
wire _1454__bF$buf3 ;
wire _1454__bF$buf4 ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _3081__bF$buf0 ;
wire _3081__bF$buf1 ;
wire _3081__bF$buf2 ;
wire _3081__bF$buf3 ;
wire _3081__bF$buf4 ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _7640_ ;
wire _7220_ ;
wire _2199_ ;
wire _8005_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _6911_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf0  ;
wire _8234_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf3  ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _7925_ ;
wire _7505_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf4  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf0  ;
wire _8043_ ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _7734_ ;
wire _7314_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _6310__bF$buf0 ;
wire _6310__bF$buf1 ;
wire _6310__bF$buf2 ;
wire _6310__bF$buf3 ;
wire _6310__bF$buf4 ;
wire _8272_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _7963_ ;
wire _7543_ ;
wire _7123_ ;
wire _8328_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf0  ;
wire _4668_ ;
wire _4248_ ;
wire [4:0] \datapath_1.a3  ;
wire _8081_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf3  ;
wire _6814_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _7772_ ;
wire _7352_ ;
wire _8137_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _7828_ ;
wire _7408_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _7581_ ;
wire _7161_ ;
wire _8366_ ;
wire _3081_ ;
wire _1814_ ;
wire _926__bF$buf0 ;
wire _4286_ ;
wire _926__bF$buf1 ;
wire _926__bF$buf2 ;
wire _926__bF$buf3 ;
wire _926__bF$buf4 ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire _7637_ ;
wire _7217_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _7390_ ;
wire _5703_ ;
wire _8175_ ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7866_ ;
wire _7446_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire _7675_ ;
wire _7255_ ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf1  ;
wire _7484_ ;
wire _7064_ ;
wire _8269_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _3869__bF$buf0 ;
wire _3869__bF$buf1 ;
wire _3869__bF$buf2 ;
wire _3869__bF$buf3 ;
wire _3869__bF$buf4 ;
wire _4821_ ;
wire _4401_ ;
wire _7293_ ;
wire _5606_ ;
wire _8078_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf1  ;
wire _190_ ;
wire _7769_ ;
wire _7349_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _7998_ ;
wire _7578_ ;
wire _7158_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf4  ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire _7387_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf1  ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _7196_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf1  ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _728__bF$buf0 ;
wire _728__bF$buf1 ;
wire _728__bF$buf2 ;
wire _728__bF$buf3 ;
wire _728__bF$buf4 ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire [31:0] _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _8002_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6250__bF$buf0 ;
wire _6250__bF$buf1 ;
wire _6250__bF$buf2 ;
wire _6085_ ;
wire _6250__bF$buf3 ;
wire _6250__bF$buf4 ;
wire _4818_ ;
wire _8231_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf0  ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _7922_ ;
wire _7502_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf1  ;
wire _4627_ ;
wire _4207_ ;
wire _7099_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf4  ;
wire _8040_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire [31:0] \datapath_1.regfile_1.regOut[19]  ;
wire _1085_ ;
wire _3084__bF$buf0 ;
wire _3084__bF$buf1 ;
wire _7731_ ;
wire _3084__bF$buf2 ;
wire _7311_ ;
wire _3084__bF$buf3 ;
wire _3084__bF$buf4 ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _7960_ ;
wire _7540_ ;
wire _7120_ ;
wire _2099_ ;
wire _8325_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf0  ;
wire _6811_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf3  ;
wire _2731_ ;
wire _2311_ ;
wire [31:0] _3936_ ;
wire _3516_ ;
wire _8134_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf4  ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf3  ;
wire _1599_ ;
wire _1179_ ;
wire _7825_ ;
wire _7405_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire _8363_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire _7634_ ;
wire _7214_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire rst_bF$buf80 ;
wire rst_bF$buf81 ;
wire rst_bF$buf82 ;
wire rst_bF$buf83 ;
wire rst_bF$buf84 ;
wire rst_bF$buf85 ;
wire rst_bF$buf86 ;
wire rst_bF$buf87 ;
wire rst_bF$buf88 ;
wire rst_bF$buf89 ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _8172_ ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire [31:0] _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7863_ ;
wire _7443_ ;
wire _7023_ ;
wire _8228_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _6714_ ;
wire _760_ ;
wire _340_ ;
wire _7919_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _7672_ ;
wire _7252_ ;
wire _8385__bF$buf0 ;
wire _8385__bF$buf1 ;
wire _8385__bF$buf2 ;
wire _8385__bF$buf3 ;
wire _8385__bF$buf4 ;
wire _8037_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _7728_ ;
wire _7308_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _7481_ ;
wire _7061_ ;
wire _8266_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _7957_ ;
wire _7537_ ;
wire _7117_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _7290_ ;
wire _5603_ ;
wire _8075_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire _7766_ ;
wire _7346_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire [31:0] _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _7995_ ;
wire _7575_ ;
wire _7155_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf1  ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _7384_ ;
wire _8169_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _7193_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf4  ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire _7669_ ;
wire _7249_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _7898_ ;
wire _7478_ ;
wire _7058_ ;
wire _2193_ ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire [31:0] _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf3  ;
wire _4815_ ;
wire _7287_ ;
wire _5773_ ;
wire _5353_ ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4624_ ;
wire _4204_ ;
wire _7096_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf1  ;
wire _5829_ ;
wire _5409_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf4  ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _8322_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf0  ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _8131_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf1  ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf0  ;
wire _1596_ ;
wire _1176_ ;
wire _7822_ ;
wire _7402_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _3087__bF$buf0 ;
wire _3087__bF$buf1 ;
wire _3087__bF$buf2 ;
wire _3087__bF$buf3 ;
wire _3087__bF$buf4 ;
wire _8360_ ;
wire _4280_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf4  ;
wire _5485_ ;
wire _5065_ ;
wire _7631_ ;
wire _7211_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire rst_bF$buf50 ;
wire rst_bF$buf51 ;
wire rst_bF$buf52 ;
wire rst_bF$buf53 ;
wire rst_bF$buf54 ;
wire rst_bF$buf55 ;
wire rst_bF$buf56 ;
wire rst_bF$buf57 ;
wire rst_bF$buf58 ;
wire rst_bF$buf59 ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _6902_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7860_ ;
wire _7440_ ;
wire _7020_ ;
wire _8225_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _7916_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf4  ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _8034_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _4200__bF$buf0 ;
wire _1499_ ;
wire _4200__bF$buf1 ;
wire _1079_ ;
wire _4200__bF$buf2 ;
wire _4200__bF$buf3 ;
wire _4200__bF$buf4 ;
wire _7725_ ;
wire _7305_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _8263_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _7954_ ;
wire _7534_ ;
wire _7114_ ;
wire _8319_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf2  ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _8072_ ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _7763_ ;
wire _7343_ ;
wire _8128_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _660_ ;
wire _240_ ;
wire _7819_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _7992_ ;
wire _7572_ ;
wire _7152_ ;
wire _8357_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _7628_ ;
wire _7208_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _7381_ ;
wire _8166_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _7857_ ;
wire _7437_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _794__bF$buf0 ;
wire _794__bF$buf1 ;
wire _794__bF$buf2 ;
wire _794__bF$buf3 ;
wire _794__bF$buf4 ;
wire _7190_ ;
wire _5923_ ;
wire _5503_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf1  ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf4  ;
wire _7666_ ;
wire _7246_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _7895_ ;
wire _7475_ ;
wire _7055_ ;
wire _2190_ ;
wire [31:0] \datapath_1.regfile_1.regOut[1]  ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf0  ;
wire _4812_ ;
wire _7284_ ;
wire _8069_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf4  ;
wire _4621_ ;
wire _4201_ ;
wire _7093_ ;
wire _5826_ ;
wire _5406_ ;
wire _8298_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf1  ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6784_ ;
wire _6364_ ;
wire _7989_ ;
wire _7569_ ;
wire _7149_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf2  ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire [31:0] \datapath_1.regfile_1.regOut[24]  ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _7798_ ;
wire _7378_ ;
wire _2093_ ;
wire _3298_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf3  ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _7187_ ;
wire _5673_ ;
wire _5253_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf1  ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf4  ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _1649_ ;
wire _1229_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf1  ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire rst_bF$buf20 ;
wire rst_bF$buf21 ;
wire rst_bF$buf22 ;
wire rst_bF$buf23 ;
wire rst_bF$buf24 ;
wire rst_bF$buf25 ;
wire rst_bF$buf26 ;
wire rst_bF$buf27 ;
wire rst_bF$buf28 ;
wire rst_bF$buf29 ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _596__bF$buf0 ;
wire _596__bF$buf1 ;
wire _596__bF$buf2 ;
wire _596__bF$buf3 ;
wire _596__bF$buf4 ;
wire _4809_ ;
wire _8222_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire [31:0] \datapath_1.mux_wd3.dout  ;
wire _1687_ ;
wire _1267_ ;
wire _7913_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf1  ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _8031_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _7722_ ;
wire _7302_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _8260_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _7951_ ;
wire _7531_ ;
wire _7111_ ;
wire _8316_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _7760_ ;
wire _7340_ ;
wire _8125_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _7816_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _4203__bF$buf0 ;
wire _4203__bF$buf1 ;
wire _4203__bF$buf2 ;
wire _4203__bF$buf3 ;
wire _4203__bF$buf4 ;
wire _8354_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _7625_ ;
wire _7205_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _6323__bF$buf0 ;
wire _6323__bF$buf1 ;
wire _6323__bF$buf2 ;
wire _8163_ ;
wire _6323__bF$buf3 ;
wire _6323__bF$buf4 ;
wire _29_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf2  ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7854_ ;
wire _7434_ ;
wire _7014_ ;
wire _8219_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf1  ;
wire _7663_ ;
wire _7243_ ;
wire _8028_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _7719_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _1388__bF$buf0 ;
wire _1388__bF$buf1 ;
wire _1388__bF$buf2 ;
wire _1388__bF$buf3 ;
wire _1388__bF$buf4 ;
wire _3639_ ;
wire _3219_ ;
wire _7892_ ;
wire _7472_ ;
wire _7052_ ;
wire _8257_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _7948_ ;
wire _7528_ ;
wire _7108_ ;
wire _2663_ ;
wire _2243_ ;
wire _4195__bF$buf0 ;
wire _4195__bF$buf1 ;
wire _4195__bF$buf2 ;
wire _4195__bF$buf3 ;
wire _4195__bF$buf4 ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _7281_ ;
wire _8066_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _7757_ ;
wire _7337_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf1  ;
wire _3677_ ;
wire _3257_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf4  ;
wire _7090_ ;
wire _5823_ ;
wire _5403_ ;
wire _8295_ ;
wire _6608_ ;
wire _1743_ ;
wire [31:0] _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _7986_ ;
wire _7566_ ;
wire _7146_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _6244__bF$buf0 ;
wire _6244__bF$buf1 ;
wire _4903_ ;
wire _6244__bF$buf2 ;
wire _6244__bF$buf3 ;
wire _6244__bF$buf4 ;
wire _7795_ ;
wire _7375_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf0  ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _7184_ ;
wire _5917_ ;
wire _8389_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf4  ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf1  ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf4  ;
wire _5726_ ;
wire _5306_ ;
wire _8198_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf2  ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _7889_ ;
wire _7469_ ;
wire _7049_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire [31:0] \datapath_1.regfile_1.regOut[14]  ;
wire _1875_ ;
wire [31:0] _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _7698_ ;
wire _7278_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _7910_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire \datapath_1.PCJump_17_bF$buf3  ;
wire _4615_ ;
wire _7087_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _68__bF$buf0 ;
wire _68__bF$buf1 ;
wire _68__bF$buf2 ;
wire _68__bF$buf3 ;
wire _68__bF$buf4 ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _6259__bF$buf0 ;
wire _6259__bF$buf1 ;
wire _6259__bF$buf2 ;
wire _6259__bF$buf3 ;
wire _6259__bF$buf4 ;
wire _2087_ ;
wire _8313_ ;
wire _4653_ ;
wire [31:0] memoryWriteData ;
wire _4233_ ;
wire [31:0] \datapath_1.regfile_1.regOut[8]  ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire _8122_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf3  ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire [31:0] _1587_ ;
wire _1167_ ;
wire _7813_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _8351_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _7622_ ;
wire _7202_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _8160_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire clk_bF$buf100 ;
wire clk_bF$buf101 ;
wire clk_bF$buf102 ;
wire clk_bF$buf103 ;
wire clk_bF$buf104 ;
wire clk_bF$buf105 ;
wire clk_bF$buf106 ;
wire _7851_ ;
wire clk_bF$buf107 ;
wire _7431_ ;
wire clk_bF$buf108 ;
wire _7011_ ;
wire clk_bF$buf109 ;
wire _8216_ ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _7907_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _7660_ ;
wire _7240_ ;
wire _8025_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _7716_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf2  ;
wire _3636_ ;
wire _3216_ ;
wire _8254_ ;
wire _1702_ ;
wire _4210__bF$buf0 ;
wire _4210__bF$buf1 ;
wire _4594_ ;
wire _4210__bF$buf2 ;
wire _4174_ ;
wire _4210__bF$buf3 ;
wire _4210__bF$buf4 ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6326__bF$buf0 ;
wire _6326__bF$buf1 ;
wire _6326__bF$buf2 ;
wire _6326__bF$buf3 ;
wire _6326__bF$buf4 ;
wire _6740_ ;
wire _6320_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf2  ;
wire _1299_ ;
wire _7945_ ;
wire _7525_ ;
wire _7105_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _8063_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _7754_ ;
wire _7334_ ;
wire _8119_ ;
wire _3674_ ;
wire _3254_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf1  ;
wire ALUSrcA ;
wire [1:0] ALUSrcB ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _8292_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _7983_ ;
wire _7563_ ;
wire _7143_ ;
wire _8348_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _880_ ;
wire _460_ ;
wire _7619_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _7792_ ;
wire _7372_ ;
wire _8157_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _7848_ ;
wire _7428_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire [3:0] _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _7181_ ;
wire _5914_ ;
wire _8386_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf1  ;
wire _1834_ ;
wire _1414_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf4  ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire _7657_ ;
wire _7237_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf1  ;
wire _5723_ ;
wire _5303_ ;
wire _8195_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf4  ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7886_ ;
wire _7466_ ;
wire _7046_ ;
wire _2181_ ;
wire _3386_ ;
wire _6247__bF$buf0 ;
wire _6247__bF$buf1 ;
wire _6247__bF$buf2 ;
wire _6247__bF$buf3 ;
wire _6247__bF$buf4 ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _7695_ ;
wire _7275_ ;
wire _3195_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire \datapath_1.PCJump_17_bF$buf0  ;
wire _4612_ ;
wire _7084_ ;
wire _5817_ ;
wire _8289_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf4  ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf2  ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _8098_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _7789_ ;
wire _7369_ ;
wire _2084_ ;
wire _8310_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _4706_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf3  ;
wire _7598_ ;
wire _7178_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf0  ;
wire _3098_ ;
wire _5664_ ;
wire _5244_ ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _7810_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _3605__bF$buf0 ;
wire _3605__bF$buf1 ;
wire _3605__bF$buf2 ;
wire _3605__bF$buf3 ;
wire _3605__bF$buf4 ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _8213_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf3  ;
wire _1678_ ;
wire _1258_ ;
wire _7904_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _8022_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _7713_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _8251_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire BranchNe ;
wire _1296_ ;
wire _7942_ ;
wire _7522_ ;
wire _7102_ ;
wire _8307_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _8060_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _7751_ ;
wire _7331_ ;
wire _8116_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _7807_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _7980_ ;
wire _7560_ ;
wire _7140_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf2  ;
wire _8345_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _7616_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _8154_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire ALUZero ;
wire _1199_ ;
wire _7845_ ;
wire _7425_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _8383_ ;
wire _1831_ ;
wire _1411_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf1  ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _7654_ ;
wire _7234_ ;
wire _8019_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _8192_ ;
wire _58_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf1  ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _7883_ ;
wire _7463_ ;
wire _7043_ ;
wire _8248_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf3  ;
wire _780_ ;
wire _360_ ;
wire _7939_ ;
wire _7519_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _7692_ ;
wire _7272_ ;
wire _8057_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf4  ;
wire _7748_ ;
wire _7328_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _7081_ ;
wire _5814_ ;
wire _8286_ ;
wire _1734_ ;
wire _1314_ ;
wire [31:0] \datapath_1.a  ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf1  ;
wire _6772_ ;
wire _6352_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf4  ;
wire _7977_ ;
wire _7557_ ;
wire _7137_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _8095_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _7786_ ;
wire _7366_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf0  ;
wire _7595_ ;
wire _7175_ ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf4  ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _8189_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _7689_ ;
wire _7269_ ;
wire _8210_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf0  ;
wire _1675_ ;
wire _1255_ ;
wire _7901_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _7498_ ;
wire _7078_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire \datapath_1.PCJump_27_bF$buf3  ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _7710_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6998_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _8304_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf3  ;
wire _8113_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _7804_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _8342_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf2  ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _7613_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _4189__bF$buf0 ;
wire _3113_ ;
wire _4189__bF$buf1 ;
wire _4189__bF$buf2 ;
wire _4189__bF$buf3 ;
wire _4189__bF$buf4 ;
wire _4738_ ;
wire _4318_ ;
wire _8151_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7842_ ;
wire _7422_ ;
wire _7002_ ;
wire _8207_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _8380_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [31:0] ALUOut ;
wire _7651_ ;
wire _7231_ ;
wire _8016_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf2  ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire _7707_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7880_ ;
wire _7460_ ;
wire _7040_ ;
wire _8245_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf2  ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf0  ;
wire _7936_ ;
wire _7516_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _8054_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf1  ;
wire _7745_ ;
wire _7325_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire [31:0] \datapath_1.alu_1.ALUInA  ;
wire _8283_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf1  ;
wire _7974_ ;
wire _7554_ ;
wire _7134_ ;
wire _8339_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _8092_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf3  ;
wire _7783_ ;
wire _7363_ ;
wire _8148_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire [31:0] _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _7839_ ;
wire _7419_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _7592_ ;
wire _7172_ ;
wire _5905_ ;
wire _8377_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire _7648_ ;
wire _7228_ ;
wire _2783_ ;
wire _2363_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf1  ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf4  ;
wire _5714_ ;
wire _8186_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _7877_ ;
wire _7457_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf4  ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _7686_ ;
wire _7266_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _7495_ ;
wire _7075_ ;
wire [31:0] \datapath_1.regfile_1.regOut[3]  ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire \datapath_1.PCJump_27_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_1_bF$buf4  ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire [1:1] PCSource ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _8089_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _8301_ ;
wire _4641_ ;
wire _4221_ ;
wire _530__bF$buf0 ;
wire _530__bF$buf1 ;
wire _530__bF$buf2 ;
wire _530__bF$buf3 ;
wire _530__bF$buf4 ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf0  ;
wire _7589_ ;
wire _7169_ ;
wire _8110_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire [2:0] ALUControl ;
wire _5655_ ;
wire _5235_ ;
wire [31:0] \datapath_1.regfile_1.regOut[26]  ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _7801_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _7398_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _7610_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf3  ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _8204_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf3  ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _4160__bF$buf0 ;
wire _4160__bF$buf1 ;
wire _5082_ ;
wire _4160__bF$buf2 ;
wire _4160__bF$buf3 ;
wire _4160__bF$buf4 ;
wire _3815_ ;
wire _6287_ ;
wire _8013_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _1850__bF$buf0 ;
wire _1850__bF$buf1 ;
wire _1850__bF$buf2 ;
wire _1850__bF$buf3 ;
wire _1850__bF$buf4 ;
wire _52_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf2  ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _7704_ ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _8242_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _7933_ ;
wire _7513_ ;
wire _198_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _8051_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _7742_ ;
wire _7322_ ;
wire _8107_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _8280_ ;
wire _2933_ ;
wire _2513_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf2  ;
wire _3718_ ;
wire _7971_ ;
wire _7551_ ;
wire _7131_ ;
wire _8336_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _7607_ ;
wire _2742_ ;
wire _2322_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf2  ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf0  ;
wire _7780_ ;
wire _7360_ ;
wire _332__bF$buf0 ;
wire _332__bF$buf1 ;
wire _332__bF$buf2 ;
wire _332__bF$buf3 ;
wire _332__bF$buf4 ;
wire _8145_ ;
wire _3280_ ;
wire _4485_ ;
wire _4223__bF$buf0 ;
wire _4223__bF$buf1 ;
wire _4065_ ;
wire _4223__bF$buf2 ;
wire _4223__bF$buf3 ;
wire _4223__bF$buf4 ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _7836_ ;
wire _7416_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _8374_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire _7645_ ;
wire _7225_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf1  ;
wire _5711_ ;
wire _8183_ ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _7874_ ;
wire _7454_ ;
wire _7034_ ;
wire _8239_ ;
wire _3794_ ;
wire _3374_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf1  ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire \datapath_1.PCJump_22_bF$buf1  ;
wire MemToReg_bF$buf0 ;
wire MemToReg_bF$buf1 ;
wire MemToReg_bF$buf2 ;
wire MemToReg_bF$buf3 ;
wire MemToReg_bF$buf4 ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _7683_ ;
wire _7263_ ;
wire _8048_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _7739_ ;
wire _7319_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _7492_ ;
wire _7072_ ;
wire _5805_ ;
wire _8277_ ;
wire _1652__bF$buf0 ;
wire _1652__bF$buf1 ;
wire _1652__bF$buf2 ;
wire _1652__bF$buf3 ;
wire _1652__bF$buf4 ;
wire _1725_ ;
wire _1305_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf4  ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf1  ;
wire _6763_ ;
wire _6343_ ;
wire _7968_ ;
wire _7548_ ;
wire _7128_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _8086_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire _7777_ ;
wire _7357_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _7586_ ;
wire _7166_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _1124__bF$buf0 ;
wire _1124__bF$buf1 ;
wire _1124__bF$buf2 ;
wire _1124__bF$buf3 ;
wire _1124__bF$buf4 ;
wire _4923_ ;
wire _4503_ ;
wire _7395_ ;
wire _5708_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf0  ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _8201_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf0  ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _3342__bF$buf0 ;
wire _3342__bF$buf1 ;
wire _3342__bF$buf2 ;
wire _5746_ ;
wire _3342__bF$buf3 ;
wire _5326_ ;
wire _3342__bF$buf4 ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _7489_ ;
wire _7069_ ;
wire _8010_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire [31:0] \datapath_1.regfile_1.regOut[16]  ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _7701_ ;
wire _386_ ;
wire clk_bF$buf90 ;
wire clk_bF$buf91 ;
wire clk_bF$buf92 ;
wire clk_bF$buf93 ;
wire clk_bF$buf94 ;
wire clk_bF$buf95 ;
wire _3621_ ;
wire clk_bF$buf96 ;
wire _3201_ ;
wire clk_bF$buf97 ;
wire clk_bF$buf98 ;
wire clk_bF$buf99 ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _7298_ ;
wire _5784_ ;
wire _5364_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf3  ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _7930_ ;
wire _7510_ ;
wire _4065__bF$buf0 ;
wire _4065__bF$buf1 ;
wire _4065__bF$buf2 ;
wire _4065__bF$buf3 ;
wire _4065__bF$buf4 ;
wire _4065__bF$buf5 ;
wire _4065__bF$buf6 ;
wire _4065__bF$buf7 ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _8104_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf2  ;
wire _8333_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _7604_ ;
wire _289_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf2  ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _8142_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _7833_ ;
wire _7413_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _8371_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _7642_ ;
wire _7222_ ;
wire _8007_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _8180_ ;
wire _46_ ;
wire _6913_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _7871_ ;
wire _7451_ ;
wire _7031_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf2  ;
wire _8236_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _7927_ ;
wire _7507_ ;
wire _2642_ ;
wire _2222_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _7680_ ;
wire _7260_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf2  ;
wire _8045_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire _4230__bF$buf0 ;
wire _4230__bF$buf1 ;
wire _4230__bF$buf2 ;
wire _4230__bF$buf3 ;
wire _4230__bF$buf4 ;
wire _7736_ ;
wire _7316_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _8274_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf1  ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _7965_ ;
wire _7545_ ;
wire _7125_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf2  ;
wire _5611_ ;
wire _8083_ ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _7774_ ;
wire _7354_ ;
wire _8139_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _7583_ ;
wire _7163_ ;
wire _8368_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire _480_ ;
wire _7639_ ;
wire _7219_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _7392_ ;
wire _5705_ ;
wire _8177_ ;
wire [31:0] \datapath_1.regfile_1.regOut[31]  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _7868_ ;
wire _7448_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire _6052_ ;
wire _7677_ ;
wire _7257_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _4151__bF$buf0 ;
wire _4151__bF$buf1 ;
wire _4151__bF$buf2 ;
wire _4151__bF$buf3 ;
wire _4151__bF$buf4 ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf3  ;
wire _7486_ ;
wire _7066_ ;
wire [31:0] _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _7295_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf0  ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf3  ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1718__bF$buf0 ;
wire _1718__bF$buf1 ;
wire _1718__bF$buf2 ;
wire _1718__bF$buf3 ;
wire _1718__bF$buf4 ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _8101_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire IRWrite ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire _7389_ ;
wire _8330_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _7601_ ;
wire _286_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf3  ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire [31:0] _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _4214__bF$buf0 ;
wire _7198_ ;
wire _4214__bF$buf1 ;
wire _4214__bF$buf2 ;
wire _4214__bF$buf3 ;
wire _4214__bF$buf4 ;
wire _5684_ ;
wire _5264_ ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _7830_ ;
wire _7410_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf3  ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _8004_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _6910_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire rst_hier0_bF$buf0 ;
wire rst_hier0_bF$buf1 ;
wire rst_hier0_bF$buf2 ;
wire rst_hier0_bF$buf3 ;
wire rst_hier0_bF$buf4 ;
wire rst_hier0_bF$buf5 ;
wire rst_hier0_bF$buf6 ;
wire rst_hier0_bF$buf7 ;
wire rst_hier0_bF$buf8 ;
wire rst_hier0_bF$buf9 ;
wire _4001__bF$buf0 ;
wire _4001__bF$buf1 ;
wire _4001__bF$buf2 ;
wire _4001__bF$buf3 ;
wire _4001__bF$buf4 ;
wire _8233_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf2  ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _7924_ ;
wire _7504_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf3  ;
wire _4629_ ;
wire _4209_ ;
wire _8042_ ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _7733_ ;
wire _7313_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _8271_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _7962_ ;
wire _7542_ ;
wire _7122_ ;
wire _8327_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _8080_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf2  ;
wire _6813_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _7771_ ;
wire _7351_ ;
wire _8136_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _7827_ ;
wire _7407_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _7580_ ;
wire _7160_ ;
wire _8365_ ;
wire _3080_ ;
wire [3:0] \control_1.next  ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire _7636_ ;
wire _7216_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _8174_ ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire ALUSrcA_bF$buf0 ;
wire _113_ ;
wire ALUSrcA_bF$buf1 ;
wire ALUSrcA_bF$buf2 ;
wire ALUSrcA_bF$buf3 ;
wire ALUSrcA_bF$buf4 ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7865_ ;
wire _7445_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire [31:0] _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _7674_ ;
wire _7254_ ;
wire _8039_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf0  ;
wire _7483_ ;
wire _7063_ ;
wire _8268_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _7959_ ;
wire _7539_ ;
wire _7119_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _7292_ ;
wire _5605_ ;
wire _8077_ ;
wire [31:0] \datapath_1.regfile_1.regOut[21]  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf0  ;
wire _7768_ ;
wire _7348_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _4154__bF$buf0 ;
wire _3900_ ;
wire _4154__bF$buf1 ;
wire _4154__bF$buf2 ;
wire _4154__bF$buf3 ;
wire _4154__bF$buf4 ;
wire _6792_ ;
wire _6372_ ;
wire _7997_ ;
wire _7577_ ;
wire _7157_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf3  ;
wire _5643_ ;
wire _5223_ ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire [31:0] _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _7386_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf0  ;
wire _4723_ ;
wire _4303_ ;
wire _7195_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf0  ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _3352__bF$buf0 ;
wire _3352__bF$buf1 ;
wire _3352__bF$buf2 ;
wire _3352__bF$buf3 ;
wire _3352__bF$buf4 ;
wire _8001_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _7289_ ;
wire _8230_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _4217__bF$buf0 ;
wire _4217__bF$buf1 ;
wire _4217__bF$buf2 ;
wire _4217__bF$buf3 ;
wire _4217__bF$buf4 ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _7921_ ;
wire _7501_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf0  ;
wire _4626_ ;
wire _4206_ ;
wire _7098_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf3  ;
wire _992__bF$buf0 ;
wire _992__bF$buf1 ;
wire _992__bF$buf2 ;
wire _992__bF$buf3 ;
wire _992__bF$buf4 ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _7730_ ;
wire _7310_ ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire _6289__bF$buf0 ;
wire _6289__bF$buf1 ;
wire _6289__bF$buf2 ;
wire _6289__bF$buf3 ;
wire _6289__bF$buf4 ;
wire _2098_ ;
wire _8324_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf2  ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _6293__bF$buf0 ;
wire _3935_ ;
wire _3515_ ;
wire _6293__bF$buf1 ;
wire _6293__bF$buf2 ;
wire _6293__bF$buf3 ;
wire _6293__bF$buf4 ;
wire _8133_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf3  ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf2  ;
wire _1598_ ;
wire _1178_ ;
wire _7824_ ;
wire _7404_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _8362_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _7633_ ;
wire _7213_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire rst_bF$buf70 ;
wire rst_bF$buf71 ;
wire rst_bF$buf72 ;
wire rst_bF$buf73 ;
wire rst_bF$buf74 ;
wire rst_bF$buf75 ;
wire rst_bF$buf76 ;
wire rst_bF$buf77 ;
wire rst_bF$buf78 ;
wire rst_bF$buf79 ;
wire [31:1] \datapath_1.regfile_1.regEn  ;
wire _4758_ ;
wire _4338_ ;
wire _8171_ ;
wire _37_ ;
wire _6904_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7862_ ;
wire _7442_ ;
wire _7022_ ;
wire _8227_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire _7918_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _7671_ ;
wire _7251_ ;
wire _8036_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _4236__bF$buf0 ;
wire _4236__bF$buf1 ;
wire _4236__bF$buf2 ;
wire _4236__bF$buf3 ;
wire _4236__bF$buf4 ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _7727_ ;
wire _7307_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _7480_ ;
wire _7060_ ;
wire _8265_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6751_ ;
wire _6331_ ;
wire _7956_ ;
wire _7536_ ;
wire _7116_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf4  ;
wire _5602_ ;
wire _8074_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire _7765_ ;
wire _7345_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _7994_ ;
wire _7574_ ;
wire _7154_ ;
wire _8359_ ;
wire _3494_ ;
wire _3074_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf0  ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _7383_ ;
wire _8168_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _7859_ ;
wire _7439_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _7192_ ;
wire _5925_ ;
wire _5505_ ;
wire [31:0] \datapath_1.regfile_1.regOut[11]  ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf3  ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire _266__bF$buf0 ;
wire _266__bF$buf1 ;
wire _266__bF$buf2 ;
wire _266__bF$buf3 ;
wire _266__bF$buf4 ;
wire _7668_ ;
wire _7248_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _7897_ ;
wire _7477_ ;
wire _7057_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf2  ;
wire _4814_ ;
wire _7286_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _4623_ ;
wire _4203_ ;
wire _7095_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf0  ;
wire [31:0] \datapath_1.regfile_1.regOut[5]  ;
wire _5828_ ;
wire _5408_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf3  ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf4  ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _1586__bF$buf0 ;
wire _1586__bF$buf1 ;
wire _1586__bF$buf2 ;
wire _1586__bF$buf3 ;
wire _2095_ ;
wire _1586__bF$buf4 ;
wire _8321_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire [31:0] \datapath_1.ALUResult  ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _7189_ ;
wire _8130_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf0  ;
wire _5675_ ;
wire _5255_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf3  ;
wire [31:0] \datapath_1.regfile_1.regOut[28]  ;
wire _1595_ ;
wire _1175_ ;
wire _7821_ ;
wire _7401_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf3  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _7630_ ;
wire _7210_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire rst_bF$buf40 ;
wire rst_bF$buf41 ;
wire rst_bF$buf42 ;
wire rst_bF$buf43 ;
wire rst_bF$buf44 ;
wire rst_bF$buf45 ;
wire rst_bF$buf46 ;
wire rst_bF$buf47 ;
wire rst_bF$buf48 ;
wire rst_bF$buf49 ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _6901_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _1058__bF$buf0 ;
wire _1058__bF$buf1 ;
wire _1058__bF$buf2 ;
wire _1058__bF$buf3 ;
wire _1058__bF$buf4 ;
wire [31:0] _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _8224_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _1689_ ;
wire _1269_ ;
wire _7915_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf3  ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _8033_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _7724_ ;
wire _7304_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _8262_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire [31:0] _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [31:0] memoryAddress ;
wire _7953_ ;
wire _7533_ ;
wire _7113_ ;
wire _8318_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf1  ;
wire _4658_ ;
wire _4238_ ;
wire _8071_ ;
wire _6804_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _7762_ ;
wire _7342_ ;
wire _8127_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire PCEn ;
wire _906_ ;
wire _6613_ ;
wire _4239__bF$buf0 ;
wire _7818_ ;
wire _4239__bF$buf1 ;
wire _4239__bF$buf2 ;
wire _4239__bF$buf3 ;
wire _4239__bF$buf4 ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire [31:0] _3738_ ;
wire _3318_ ;
wire _7991_ ;
wire _7571_ ;
wire _7151_ ;
wire _8356_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _7627_ ;
wire _7207_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _7380_ ;
wire _8165_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf4  ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7856_ ;
wire _7436_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire [31:0] _333_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf0  ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf3  ;
wire _7665_ ;
wire _7245_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire [31:0] _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _7894_ ;
wire _7474_ ;
wire _7054_ ;
wire _8259_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _7283_ ;
wire _8068_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire [31:8] \datapath_1.PCJump  ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _7759_ ;
wire _7339_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf3  ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _7092_ ;
wire _5825_ ;
wire _5405_ ;
wire _8297_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf0  ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _7988_ ;
wire _7568_ ;
wire _7148_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf1  ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire [31:0] _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _7797_ ;
wire _7377_ ;
wire _2092_ ;
wire _3297_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf2  ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _7186_ ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf0  ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf3  ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf4  ;
wire _1648_ ;
wire _1228_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf0  ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire rst_bF$buf10 ;
wire rst_bF$buf11 ;
wire rst_bF$buf12 ;
wire rst_bF$buf13 ;
wire rst_bF$buf14 ;
wire rst_bF$buf15 ;
wire rst_bF$buf16 ;
wire rst_bF$buf17 ;
wire rst_bF$buf18 ;
wire rst_bF$buf19 ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _4808_ ;
wire _8221_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _7912_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf0  ;
wire [31:0] _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _7089_ ;
wire _8030_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire [31:0] \datapath_1.regfile_1.regOut[18]  ;
wire _1495_ ;
wire _1075_ ;
wire _7721_ ;
wire _7301_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _7950_ ;
wire _7530_ ;
wire _7110_ ;
wire _2089_ ;
wire _8315_ ;
wire [31:0] _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _4183__bF$buf0 ;
wire _4183__bF$buf1 ;
wire _4183__bF$buf2 ;
wire _4183__bF$buf3 ;
wire _4183__bF$buf4 ;
wire _6801_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _8124_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _1589_ ;
wire _1169_ ;
wire _7815_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _8353_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _7624_ ;
wire _7204_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _8162_ ;
wire _28_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf1  ;
wire _1610_ ;
wire _6232__bF$buf0 ;
wire _6232__bF$buf1 ;
wire _6232__bF$buf2 ;
wire _6232__bF$buf3 ;
wire _6232__bF$buf4 ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire [27:0] \datapath_1.mux_iord.din0  ;
wire _7853_ ;
wire _7433_ ;
wire _7013_ ;
wire _8218_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _6704_ ;
wire _750_ ;
wire _330_ ;
wire _7909_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf0  ;
wire _3829_ ;
wire _3409_ ;
wire _7662_ ;
wire _7242_ ;
wire _8027_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _7718_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf4  ;
wire _3638_ ;
wire _3218_ ;
wire _7891_ ;
wire _7471_ ;
wire _7051_ ;
wire _8256_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf4  ;
wire _7947_ ;
wire _7527_ ;
wire _7107_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _7280_ ;
wire _8065_ ;
wire _3803__bF$buf0 ;
wire _3803__bF$buf1 ;
wire _3803__bF$buf2 ;
wire _3803__bF$buf3 ;
wire _3803__bF$buf4 ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _7756_ ;
wire _7336_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf0  ;
wire _3676_ ;
wire _3256_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf3  ;
wire _5822_ ;
wire _5402_ ;
wire _8294_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _7985_ ;
wire _7565_ ;
wire _7145_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _7794_ ;
wire _7374_ ;
wire _8159_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _7183_ ;
wire _5916_ ;
wire _8388_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf3  ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf0  ;
wire _7659_ ;
wire _7239_ ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf3  ;
wire _5725_ ;
wire _5305_ ;
wire _8197_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf1  ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _4167__bF$buf0 ;
wire _4167__bF$buf1 ;
wire _4167__bF$buf2 ;
wire _4167__bF$buf3 ;
wire _4167__bF$buf4 ;
wire _6683_ ;
wire _6263_ ;
wire _7888_ ;
wire _7468_ ;
wire _7048_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire _7697_ ;
wire _7277_ ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire \datapath_1.PCJump_17_bF$buf2  ;
wire _4614_ ;
wire _7086_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf4  ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire _8312_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire _8121_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf2  ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _7812_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _8350_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _7621_ ;
wire _7201_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7850_ ;
wire _7430_ ;
wire _7010_ ;
wire _8215_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _7906_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _8024_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _7715_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf1  ;
wire _3635_ ;
wire _3215_ ;
wire _8253_ ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf1  ;
wire _1298_ ;
wire _7944_ ;
wire _7524_ ;
wire _7104_ ;
wire _8309_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _8062_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _7753_ ;
wire _7333_ ;
wire _8118_ ;
wire _3673_ ;
wire _3253_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf0  ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _8291_ ;
wire _6604_ ;
wire _650_ ;
wire _230_ ;
wire _7809_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _7982_ ;
wire _7562_ ;
wire _7142_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf4  ;
wire _8347_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _7618_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _7791_ ;
wire _7371_ ;
wire _8156_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _7847_ ;
wire _7427_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _7180_ ;
wire _5913_ ;
wire _8385_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf0  ;
wire _1833_ ;
wire _1413_ ;
wire IorD_bF$buf0 ;
wire IorD_bF$buf1 ;
wire IorD_bF$buf2 ;
wire IorD_bF$buf3 ;
wire IorD_bF$buf4 ;
wire \datapath_1.mux_wd3.dout_16_bF$buf3  ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire _7656_ ;
wire _7236_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf0  ;
wire _5722_ ;
wire _5302_ ;
wire _8194_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf3  ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _7885_ ;
wire _7465_ ;
wire _7045_ ;
wire _2180_ ;
wire [31:0] \datapath_1.regfile_1.regOut[0]  ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6302__bF$buf0 ;
wire _6302__bF$buf1 ;
wire _6302__bF$buf2 ;
wire _6302__bF$buf3 ;
wire _6302__bF$buf4 ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _7694_ ;
wire _7274_ ;
wire _8059_ ;
wire _3194_ ;
wire [31:0] \datapath_1.rd2  ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _7083_ ;
wire _5816_ ;
wire _8288_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf3  ;
wire _6774_ ;
wire _6354_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf1  ;
wire _7979_ ;
wire _7559_ ;
wire _7139_ ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _8097_ ;
wire [31:0] \datapath_1.regfile_1.regOut[23]  ;
wire _1965_ ;
wire _1545_ ;
wire [31:0] _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire [31:0] memoryOutData ;
wire _7788_ ;
wire _7368_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire [1:0] ALUOp ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _4705_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf2  ;
wire _7597_ ;
wire _7177_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _6317__bF$buf0 ;
wire _6317__bF$buf1 ;
wire _6317__bF$buf2 ;
wire _6317__bF$buf3 ;
wire _6317__bF$buf4 ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;
wire _8212_ ;

OR2X2 _11689_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .B(_1718__bF$buf0),
    .Y(_1658_)
);

DFFSR _11269_ (
    .CLK(clk_bF$buf48),
    .D(_1389_[7]),
    .Q(\datapath_1.regfile_1.regOut[22] [7]),
    .R(rst_bF$buf48),
    .S(vdd)
);

FILL FILL_1__13352_ (
);

AND2X2 _17915_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_6833_)
);

OR2X2 _12630_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(_2194_),
    .Y(_2195_)
);

FILL FILL_0__12345_ (
);

OR2X2 _12210_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_1925_)
);

FILL FILL505400x9880 (
);

FILL FILL434720x227240 (
);

OR2X2 _9837_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_723_)
);

OR2X2 _9417_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_503_)
);

FILL FILL_1__8794_ (
);

FILL FILL42560x281580 (
);

FILL FILL_1__14557_ (
);

OR2X2 _13835_ (
    .A(\datapath_1.a [6]),
    .B(_3342__bF$buf0),
    .Y(_3290_)
);

NAND3X1 _13415_ (
    .A(_2383_),
    .B(ALUControl[1]),
    .C(_2177_),
    .Y(_2950_)
);

FILL FILL356440x330980 (
);

FILL FILL114760x14820 (
);

DFFSR _9590_ (
    .CLK(clk_bF$buf66),
    .D(_531_[5]),
    .Q(\datapath_1.regfile_1.regOut[9] [5]),
    .R(rst_bF$buf80),
    .S(vdd)
);

AND2X2 _9170_ (
    .A(_378_),
    .B(_377_),
    .Y(_333_[22])
);

FILL FILL82080x281580 (
);

FILL FILL117800x79040 (
);

FILL FILL301720x79040 (
);

FILL FILL_0__10831_ (
);

FILL FILL_0__10411_ (
);

OR2X2 _18873_ (
    .A(_7774_),
    .B(_7775_),
    .Y(_7776_)
);

FILL FILL_0__18588_ (
);

FILL FILL_0__18168_ (
);

FILL FILL_0_BUFX2_insert901 (
);

OR2X2 _18453_ (
    .A(_7360_),
    .B(_7361_),
    .Y(_7362_)
);

AND2X2 _18033_ (
    .A(_6293__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_6949_)
);

FILL FILL_0_BUFX2_insert903 (
);

FILL FILL_0_BUFX2_insert904 (
);

FILL FILL_0_BUFX2_insert905 (
);

FILL FILL_0_BUFX2_insert906 (
);

FILL FILL_0_BUFX2_insert907 (
);

FILL FILL_0_BUFX2_insert909 (
);

FILL FILL104880x316160 (
);

FILL FILL_0__11616_ (
);

OR2X2 _11901_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_1779_)
);

FILL FILL340480x133380 (
);

AND2X2 _19238_ (
    .A(_6244__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_8135_)
);

FILL FILL380000x242060 (
);

OR2X2 _14793_ (
    .A(\datapath_1.rd2 [12]),
    .B(_3935__bF$buf1),
    .Y(_3895_)
);

OR2X2 _14373_ (
    .A(memoryOutData[1]),
    .B(_3737__bF$buf1),
    .Y(_3675_)
);

FILL FILL413440x54340 (
);

FILL FILL318440x113620 (
);

FILL FILL312360x266760 (
);

AND2X2 _15998_ (
    .A(_4239__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_4944_)
);

AND2X2 _15578_ (
    .A(_4183__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_4531_)
);

NOR2X1 _15158_ (
    .A(_4120_),
    .B(\datapath_1.a3 [1]),
    .Y(_4121_)
);

OR2X2 _10293_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_947_)
);

FILL FILL229520x276640 (
);

FILL FILL_0__16234_ (
);

FILL FILL193040x316160 (
);

FILL FILL280440x321100 (
);

AND2X2 _8861_ (
    .A(_212_),
    .B(_211_),
    .Y(_201_[5])
);

BUFX2 _8441_ (
    .A(_2_[17]),
    .Y(memoryWriteData[17])
);

FILL FILL16720x64220 (
);

AND2X2 _11498_ (
    .A(_1570_),
    .B(_1569_),
    .Y(_1521_[24])
);

FILL FILL_1__18446_ (
);

AND2X2 _11078_ (
    .A(_1350_),
    .B(_1349_),
    .Y(_1323_[13])
);

FILL FILL_0__17439_ (
);

AND2X2 _17724_ (
    .A(_6321__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_6645_)
);

FILL FILL_0__17019_ (
);

AND2X2 _17304_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_6230_)
);

FILL FILL_0__12994_ (
);

FILL FILL_0__12574_ (
);

FILL FILL125400x83980 (
);

FILL FILL_0__12154_ (
);

OR2X2 _9646_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .B(_662__bF$buf1),
    .Y(_616_)
);

DFFSR _9226_ (
    .CLK(clk_bF$buf72),
    .D(_333_[28]),
    .Q(\datapath_1.regfile_1.regOut[6] [28]),
    .R(rst_bF$buf32),
    .S(vdd)
);

FILL FILL61560x261820 (
);

AND2X2 _18929_ (
    .A(_6262__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_7831_)
);

OR2X2 _18509_ (
    .A(_7416_),
    .B(_7417_),
    .Y(_7418_)
);

FILL FILL365560x172900 (
);

FILL FILL_0__13779_ (
);

FILL FILL_0__13359_ (
);

AND2X2 _13644_ (
    .A(_3089__bF$buf2),
    .B(gnd),
    .Y(_3132_)
);

NOR3X1 _13224_ (
    .A(_2498_),
    .B(_2770_),
    .C(_2244_),
    .Y(_2771_)
);

FILL FILL_0__14720_ (
);

FILL FILL304760x281580 (
);

FILL FILL295640x177840 (
);

FILL FILL_0__17192_ (
);

OR2X2 _14849_ (
    .A(vdd),
    .B(_2_[31]),
    .Y(_3932_)
);

OR2X2 _14429_ (
    .A(vdd),
    .B(\datapath_1.Data [20]),
    .Y(_3712_)
);

AND2X2 _14009_ (
    .A(_3344__bF$buf3),
    .B(gnd),
    .Y(_3427_)
);

FILL FILL_1__16512_ (
);

FILL FILL_0_CLKBUF1_insert131 (
);

FILL FILL_0_CLKBUF1_insert132 (
);

FILL FILL_0_CLKBUF1_insert133 (
);

FILL FILL_0_CLKBUF1_insert134 (
);

FILL FILL_0_CLKBUF1_insert135 (
);

FILL FILL_0_CLKBUF1_insert137 (
);

FILL FILL_0__10220_ (
);

FILL FILL_0_CLKBUF1_insert139 (
);

FILL FILL272080x242060 (
);

OR2X2 _18682_ (
    .A(_7587_),
    .B(_7586_),
    .Y(_7588_)
);

FILL FILL_0__18397_ (
);

OR2X2 _18262_ (
    .A(_7170_),
    .B(_7173_),
    .Y(_7174_)
);

FILL FILL208240x296400 (
);

FILL FILL54720x306280 (
);

FILL FILL_0__8498_ (
);

DFFSR _10769_ (
    .CLK(clk_bF$buf82),
    .D(_1125_[23]),
    .Q(\datapath_1.regfile_1.regOut[18] [23]),
    .R(rst_bF$buf94),
    .S(vdd)
);

AND2X2 _10349_ (
    .A(_984_),
    .B(_983_),
    .Y(_927_[28])
);

FILL FILL_1__12852_ (
);

FILL FILL358720x217360 (
);

FILL FILL_1__12012_ (
);

FILL FILL_0__11845_ (
);

OR2X2 _11710_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .B(_1718__bF$buf0),
    .Y(_1672_)
);

OR2X2 _19467_ (
    .A(gnd),
    .B(_8385__bF$buf1),
    .Y(_8347_)
);

NOR2X1 _19047_ (
    .A(_6310__bF$buf4),
    .B(_7946_),
    .Y(_7947_)
);

OR2X2 _14182_ (
    .A(MemToReg_bF$buf0),
    .B(ALUOut[13]),
    .Y(_3566_)
);

OR2X2 _8917_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .B(_266__bF$buf1),
    .Y(_250_)
);

FILL FILL136800x49400 (
);

FILL FILL_1__13217_ (
);

FILL FILL471200x261820 (
);

OR2X2 _12915_ (
    .A(_2479_),
    .B(_2475_),
    .Y(_2480_)
);

FILL FILL_1_BUFX2_insert456 (
);

FILL FILL_1_BUFX2_insert458 (
);

AND2X2 _15387_ (
    .A(_4146__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_4343_)
);

FILL FILL187720x286520 (
);

FILL FILL_0__16883_ (
);

FILL FILL_0__16463_ (
);

FILL FILL_0__16043_ (
);

FILL FILL187720x83980 (
);

FILL FILL371640x83980 (
);

FILL FILL215080x9880 (
);

FILL FILL101840x350740 (
);

FILL FILL274360x197600 (
);

OR2X2 _8670_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_125_)
);

FILL FILL119320x247000 (
);

FILL FILL_0__17668_ (
);

OR2X2 _17953_ (
    .A(_6869_),
    .B(_6868_),
    .Y(_6870_)
);

AND2X2 _17533_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_6457_)
);

OR2X2 _17113_ (
    .A(_6026_),
    .B(_6041_),
    .Y(_6042_)
);

FILL FILL423320x182780 (
);

FILL FILL_0__12383_ (
);

FILL FILL294120x0 (
);

FILL FILL234080x9880 (
);

OR2X2 _9875_ (
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .Y(_793_)
);

AND2X2 _9455_ (
    .A(_528_),
    .B(_527_),
    .Y(_465_[31])
);

AND2X2 _9035_ (
    .A(_308_),
    .B(_307_),
    .Y(_267_[20])
);

FILL FILL_1__11703_ (
);

FILL FILL_1__14175_ (
);

OR2X2 _18738_ (
    .A(_7639_),
    .B(_7642_),
    .Y(_7643_)
);

OR2X2 _18318_ (
    .A(_7198_),
    .B(_7229_),
    .Y(_7230_)
);

OR2X2 _13873_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [19]),
    .Y(_3315_)
);

FILL FILL_0__13168_ (
);

AND2X2 _13453_ (
    .A(_2984_),
    .B(_2985_),
    .Y(_2986_)
);

AOI22X1 _13033_ (
    .A(_2590_),
    .B(_2548_),
    .C(_2477_),
    .D(_2504_),
    .Y(_2591_)
);

FILL FILL171760x49400 (
);

FILL FILL181640x227240 (
);

FILL FILL_1__9197_ (
);

FILL FILL323760x261820 (
);

FILL FILL_0__9915_ (
);

FILL FILL256880x4940 (
);

FILL FILL373160x316160 (
);

OR2X2 _14658_ (
    .A(\datapath_1.rd1 [10]),
    .B(_3869__bF$buf3),
    .Y(_3825_)
);

AND2X2 _14238_ (
    .A(_3603_),
    .B(_3602_),
    .Y(\datapath_1.mux_wd3.dout [31])
);

FILL FILL_1__16741_ (
);

FILL FILL_0__15734_ (
);

FILL FILL_0__15314_ (
);

OR2X2 _18491_ (
    .A(_7398_),
    .B(_7399_),
    .Y(_7400_)
);

OR2X2 _18071_ (
    .A(_6984_),
    .B(_6985_),
    .Y(_6986_)
);

FILL FILL266760x74100 (
);

OR2X2 _10998_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_1317_)
);

OR2X2 _10578_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_1097_)
);

OR2X2 _10158_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_877_)
);

FILL FILL_0__16939_ (
);

FILL FILL_0__16519_ (
);

AND2X2 _16804_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_5738_)
);

FILL FILL_0__11234_ (
);

OR2X2 _19276_ (
    .A(_8165_),
    .B(_8172_),
    .Y(_8173_)
);

AND2X2 _8726_ (
    .A(_142_),
    .B(_141_),
    .Y(_135_[3])
);

FILL FILL_0__12859_ (
);

OR2X2 _12724_ (
    .A(_2280_),
    .B(_2288_),
    .Y(_2289_)
);

DFFSR _12304_ (
    .CLK(clk_bF$buf76),
    .D(_1917_[10]),
    .Q(\datapath_1.regfile_1.regOut[30] [10]),
    .R(rst_bF$buf110),
    .S(vdd)
);

FILL FILL329080x158080 (
);

FILL FILL416480x163020 (
);

NOR3X1 _15196_ (
    .A(_4150_),
    .B(_4144_),
    .C(_4153_),
    .Y(_4154_)
);

FILL FILL_0__13800_ (
);

FILL FILL_1__8888_ (
);

FILL FILL_0__16692_ (
);

FILL FILL_0__16272_ (
);

FILL FILL481080x345800 (
);

FILL FILL329840x118560 (
);

AND2X2 _13929_ (
    .A(_3352__bF$buf2),
    .B(gnd),
    .Y(_3359_)
);

AND2X2 _13509_ (
    .A(_3027_),
    .B(_3026_),
    .Y(_1_[6])
);

FILL FILL475000x301340 (
);

FILL FILL_1__18484_ (
);

FILL FILL_1__18064_ (
);

FILL FILL209000x232180 (
);

OR2X2 _17762_ (
    .A(_6680_),
    .B(_6681_),
    .Y(_6682_)
);

FILL FILL_0__17057_ (
);

OR2X2 _17342_ (
    .A(_6253_),
    .B(_6267_),
    .Y(_6268_)
);

FILL FILL439280x113620 (
);

OR2X2 _9684_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_641_)
);

OR2X2 _9264_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_421_)
);

FILL FILL_1_CLKBUF1_insert162 (
);

FILL FILL372400x167960 (
);

FILL FILL_1__11512_ (
);

FILL FILL_1_CLKBUF1_insert164 (
);

FILL FILL_1_CLKBUF1_insert166 (
);

FILL FILL_0__10925_ (
);

FILL FILL46360x365560 (
);

OR2X2 _18967_ (
    .A(_7852_),
    .B(_7868_),
    .Y(_7869_)
);

FILL FILL177080x256880 (
);

AND2X2 _18547_ (
    .A(_6259__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_7455_)
);

AND2X2 _18127_ (
    .A(_6312__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .Y(_7041_)
);

FILL FILL_0__13397_ (
);

AND2X2 _13682_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[13]),
    .Y(_3164_)
);

AND2X2 _13262_ (
    .A(_2806_),
    .B(_2795_),
    .Y(_2807_)
);

FILL FILL95760x163020 (
);

FILL FILL_0__19203_ (
);

FILL FILL_1__12717_ (
);

FILL FILL367840x286520 (
);

FILL FILL_0__9304_ (
);

FILL FILL_1__15189_ (
);

FILL FILL505400x202540 (
);

AND2X2 _14887_ (
    .A(_3937_),
    .B(_4000_),
    .Y(_3936_[0])
);

DFFSR _14467_ (
    .CLK(clk_bF$buf65),
    .D(_3672_[2]),
    .Q(\datapath_1.Data [2]),
    .R(rst_bF$buf26),
    .S(vdd)
);

AND2X2 _14047_ (
    .A(_3350__bF$buf4),
    .B(_2_[18]),
    .Y(_3460_)
);

FILL FILL121600x59280 (
);

FILL FILL_0__15963_ (
);

FILL FILL238640x9880 (
);

FILL FILL_0__15543_ (
);

FILL FILL353400x113620 (
);

DFFSR _10387_ (
    .CLK(clk_bF$buf61),
    .D(_927_[28]),
    .Q(\datapath_1.regfile_1.regOut[15] [28]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL_1__12470_ (
);

FILL FILL_0__16748_ (
);

AND2X2 _16613_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_5550_)
);

FILL FILL257640x9880 (
);

FILL FILL484120x232180 (
);

FILL FILL247000x266760 (
);

FILL FILL_0__11463_ (
);

FILL FILL_0__11043_ (
);

AND2X2 _19085_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_7985_)
);

DFFSR _8955_ (
    .CLK(clk_bF$buf90),
    .D(_201_[15]),
    .Q(\datapath_1.regfile_1.regOut[4] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL123880x54340 (
);

OR2X2 _8535_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_55_)
);

FILL FILL_1__13675_ (
);

AND2X2 _17818_ (
    .A(_6315__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [7]),
    .Y(_6737_)
);

FILL FILL276640x9880 (
);

FILL FILL_0__12668_ (
);

NAND2X1 _12953_ (
    .A(_2379__bF$buf3),
    .B(_2353_),
    .Y(_2516_)
);

AND2X2 _12533_ (
    .A(_2122_),
    .B(_2110_),
    .Y(_2123_)
);

AND2X2 _12113_ (
    .A(_1880_),
    .B(_1879_),
    .Y(_1851_[14])
);

FILL FILL_1_BUFX2_insert835 (
);

FILL FILL_1_BUFX2_insert837 (
);

FILL FILL_1_BUFX2_insert839 (
);

FILL FILL384560x311220 (
);

FILL FILL329080x296400 (
);

FILL FILL259920x4940 (
);

AND2X2 _13738_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[21]),
    .Y(_3212_)
);

OR2X2 _13318_ (
    .A(_2849_),
    .B(_2858_),
    .Y(_2859_)
);

FILL FILL372400x98800 (
);

BUFX2 BUFX2_insert500 (
    .A(_4160_),
    .Y(_4160__bF$buf0)
);

BUFX2 BUFX2_insert501 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf4 )
);

BUFX2 BUFX2_insert502 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf3 )
);

BUFX2 BUFX2_insert503 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf2 )
);

BUFX2 BUFX2_insert504 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf1 )
);

OR2X2 _17991_ (
    .A(_6900_),
    .B(_6907_),
    .Y(_6908_)
);

AND2X2 _17571_ (
    .A(_6238__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_6494_)
);

BUFX2 BUFX2_insert505 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf0 )
);

FILL FILL_0__17286_ (
);

BUFX2 BUFX2_insert506 (
    .A(_4195_),
    .Y(_4195__bF$buf4)
);

AND2X2 _17151_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_6079_)
);

BUFX2 BUFX2_insert507 (
    .A(_4195_),
    .Y(_4195__bF$buf3)
);

BUFX2 BUFX2_insert508 (
    .A(_4195_),
    .Y(_4195__bF$buf2)
);

BUFX2 BUFX2_insert509 (
    .A(_4195_),
    .Y(_4195__bF$buf1)
);

FILL FILL118560x108680 (
);

OR2X2 _9493_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .B(_596__bF$buf2),
    .Y(_534_)
);

FILL FILL_1__16606_ (
);

DFFSR _9073_ (
    .CLK(clk_bF$buf82),
    .D(_267_[4]),
    .Q(\datapath_1.regfile_1.regOut[5] [4]),
    .R(rst_bF$buf94),
    .S(vdd)
);

FILL FILL_1__11321_ (
);

FILL FILL_0__10734_ (
);

FILL FILL_0__10314_ (
);

FILL FILL_0_BUFX2_insert21 (
);

AND2X2 _18776_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_7680_)
);

FILL FILL_0_BUFX2_insert22 (
);

FILL FILL_0_BUFX2_insert23 (
);

AND2X2 _18356_ (
    .A(_6216__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_7267_)
);

FILL FILL_0_BUFX2_insert24 (
);

FILL FILL_0_BUFX2_insert25 (
);

FILL FILL_0_BUFX2_insert27 (
);

AND2X2 _13491_ (
    .A(_3015_),
    .B(_3078_),
    .Y(_1_[0])
);

AOI21X1 _13071_ (
    .A(_2260_),
    .B(_2261_),
    .C(_2501_),
    .Y(_2627_)
);

FILL FILL_0_BUFX2_insert29 (
);

FILL FILL236360x326040 (
);

FILL FILL170240x182780 (
);

FILL FILL_0__19432_ (
);

FILL FILL183920x59280 (
);

FILL FILL503880x88920 (
);

FILL FILL222680x350740 (
);

FILL FILL_0__11519_ (
);

FILL FILL_0__9113_ (
);

DFFSR _11804_ (
    .CLK(clk_bF$buf109),
    .D(_1653_[26]),
    .Q(\datapath_1.regfile_1.regOut[26] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL203680x187720 (
);

FILL FILL184680x143260 (
);

FILL FILL243200x296400 (
);

FILL FILL152760x355680 (
);

OR2X2 _14696_ (
    .A(vdd),
    .B(\datapath_1.a [23]),
    .Y(_3850_)
);

OR2X2 _14276_ (
    .A(vdd),
    .B(ALUOut[12]),
    .Y(_3630_)
);

FILL FILL311600x39520 (
);

FILL FILL_0__15352_ (
);

FILL FILL_1__17564_ (
);

AND2X2 _10196_ (
    .A(_902_),
    .B(_901_),
    .Y(_861_[20])
);

FILL FILL34960x276640 (
);

FILL FILL357960x350740 (
);

FILL FILL231800x54340 (
);

FILL FILL_0__16557_ (
);

AND2X2 _16842_ (
    .A(_4160__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_5775_)
);

FILL FILL_0__16137_ (
);

OR2X2 _16422_ (
    .A(_5360_),
    .B(_5361_),
    .Y(_5362_)
);

AND2X2 _16002_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_4948_)
);

FILL FILL_0__11692_ (
);

OR2X2 _8764_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .B(_200__bF$buf0),
    .Y(_168_)
);

AND2X2 _17627_ (
    .A(_6321__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_6549_)
);

OR2X2 _17207_ (
    .A(_6134_),
    .B(_6127_),
    .Y(_6135_)
);

FILL FILL_0__12897_ (
);

NAND2X1 _12762_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2327_)
);

OR2X2 _12342_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_1993_)
);

FILL FILL_0__18703_ (
);

OR2X2 _9969_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_791_)
);

OR2X2 _9549_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_571_)
);

OR2X2 _9129_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_351_)
);

FILL FILL483360x34580 (
);

FILL FILL6840x54340 (
);

FILL FILL_1__14689_ (
);

FILL FILL_0_BUFX2_insert490 (
);

FILL FILL_0_BUFX2_insert492 (
);

AND2X2 _13967_ (
    .A(_3344__bF$buf0),
    .B(gnd),
    .Y(_3391_)
);

FILL FILL_0_BUFX2_insert494 (
);

OR2X2 _13547_ (
    .A(ALUOut[19]),
    .B(_3079__bF$buf4),
    .Y(_3053_)
);

OR2X2 _13127_ (
    .A(_2277_),
    .B(_2679_),
    .Y(_2680_)
);

FILL FILL_0_BUFX2_insert496 (
);

FILL FILL_0_BUFX2_insert498 (
);

FILL FILL_0_BUFX2_insert499 (
);

FILL FILL_1__15630_ (
);

FILL FILL_1__15210_ (
);

FILL FILL_0__14203_ (
);

FILL FILL162640x39520 (
);

OR2X2 _17380_ (
    .A(_6305_),
    .B(_6292_),
    .Y(_6306_)
);

FILL FILL337440x49400 (
);

FILL FILL271320x256880 (
);

FILL FILL294880x242060 (
);

FILL FILL_0__15828_ (
);

FILL FILL_0__15408_ (
);

FILL FILL_0__10963_ (
);

FILL FILL_0__10543_ (
);

FILL FILL72200x247000 (
);

AND2X2 _18585_ (
    .A(_6312__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_7492_)
);

OR2X2 _18165_ (
    .A(_7077_),
    .B(_7078_),
    .Y(_7079_)
);

FILL FILL336680x370500 (
);

FILL FILL_0__11748_ (
);

OR2X2 _11613_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_1627_)
);

FILL FILL_0__11328_ (
);

FILL FILL166440x39520 (
);

OR2X2 _14085_ (
    .A(_3492_),
    .B(_3489_),
    .Y(\datapath_1.alu_1.ALUInB [23])
);

FILL FILL_0__15581_ (
);

FILL FILL_0__15161_ (
);

NOR2X1 _12818_ (
    .A(_2154_),
    .B(_2378_),
    .Y(_2383_)
);

FILL FILL468920x64220 (
);

FILL FILL421040x207480 (
);

FILL FILL408120x88920 (
);

FILL FILL_0__16786_ (
);

AND2X2 _16651_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_5587_)
);

FILL FILL445360x64220 (
);

OR2X2 _16231_ (
    .A(_5173_),
    .B(_5170_),
    .Y(_5174_)
);

FILL FILL_0__11081_ (
);

AND2X2 _8993_ (
    .A(_280_),
    .B(_279_),
    .Y(_267_[6])
);

DFFSR _8573_ (
    .CLK(clk_bF$buf46),
    .D(_3_[20]),
    .Q(\datapath_1.regfile_1.regOut[1] [20]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL_1__10401_ (
);

FILL FILL_1__18578_ (
);

FILL FILL_1__13293_ (
);

OR2X2 _17856_ (
    .A(_6773_),
    .B(_6774_),
    .Y(_6775_)
);

AND2X2 _17436_ (
    .A(_6250__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_6361_)
);

OR2X2 _17016_ (
    .A(_5946_),
    .B(_5931_),
    .Y(_5947_)
);

NAND2X1 _12991_ (
    .A(_2551_),
    .B(_2549_),
    .Y(_2552_)
);

OR2X2 _12571_ (
    .A(\control_1.reg_state.dout [0]),
    .B(vdd),
    .Y(_2144_)
);

FILL FILL_0__12286_ (
);

OR2X2 _12151_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .B(_1916__bF$buf2),
    .Y(_1906_)
);

FILL FILL177840x326040 (
);

FILL FILL_0__18512_ (
);

FILL FILL88920x24700 (
);

OR2X2 _9778_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .B(_728__bF$buf2),
    .Y(_684_)
);

DFFSR _9358_ (
    .CLK(clk_bF$buf95),
    .D(_399_[31]),
    .Q(\datapath_1.regfile_1.regOut[7] [31]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL3800x138320 (
);

FILL FILL_0__8613_ (
);

FILL FILL_1__14498_ (
);

FILL FILL364800x0 (
);

AND2X2 _13776_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [26]),
    .Y(_3245_)
);

OAI21X1 _13356_ (
    .A(_2893_),
    .B(_2376__bF$buf0),
    .C(_2894_),
    .Y(_2895_)
);

FILL FILL3040x365560 (
);

FILL FILL_0__14432_ (
);

FILL FILL485640x182780 (
);

FILL FILL_0__14012_ (
);

FILL FILL81320x365560 (
);

FILL FILL_0__9818_ (
);

FILL FILL313120x316160 (
);

FILL FILL400520x321100 (
);

FILL FILL104880x202540 (
);

FILL FILL_0__15637_ (
);

OR2X2 _15922_ (
    .A(_4868_),
    .B(_4869_),
    .Y(_4870_)
);

AND2X2 _15502_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_4456_)
);

FILL FILL_0__15217_ (
);

FILL FILL85120x286520 (
);

FILL FILL_0__10352_ (
);

FILL FILL399760x237120 (
);

AND2X2 _18394_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_7304_)
);

FILL FILL389120x197600 (
);

FILL FILL268280x345800 (
);

FILL FILL_0__19470_ (
);

FILL FILL_0__19050_ (
);

FILL FILL_1__17429_ (
);

FILL FILL_1__12564_ (
);

AND2X2 _16707_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_5642_)
);

FILL FILL_0__11977_ (
);

FILL FILL_0__9151_ (
);

OR2X2 _11842_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_1784__bF$buf1),
    .Y(_1740_)
);

DFFSR _11422_ (
    .CLK(clk_bF$buf100),
    .D(_1455_[31]),
    .Q(\datapath_1.regfile_1.regOut[23] [31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

OR2X2 _11002_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .B(_1322__bF$buf2),
    .Y(_1320_)
);

OR2X2 _19179_ (
    .A(_8073_),
    .B(_8076_),
    .Y(_8077_)
);

OR2X2 _8629_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .B(_134__bF$buf1),
    .Y(_98_)
);

FILL FILL_0__15390_ (
);

FILL FILL_1__13769_ (
);

OR2X2 _12627_ (
    .A(_2188_),
    .B(_2191_),
    .Y(_2192_)
);

OR2X2 _12207_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_1923_)
);

FILL FILL_1__14710_ (
);

FILL FILL142880x370500 (
);

OAI21X1 _15099_ (
    .A(_4079_),
    .B(_4081_),
    .C(_4017_),
    .Y(_4082_)
);

FILL FILL_0__13703_ (
);

FILL FILL256880x118560 (
);

FILL FILL_1__17182_ (
);

AND2X2 _16880_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_5813_)
);

FILL FILL_0__16175_ (
);

OR2X2 _16460_ (
    .A(_5398_),
    .B(_5397_),
    .Y(_5399_)
);

OR2X2 _16040_ (
    .A(_4978_),
    .B(_4985_),
    .Y(_4986_)
);

FILL FILL76000x93860 (
);

FILL FILL282720x251940 (
);

FILL FILL_1__9312_ (
);

FILL FILL117800x163020 (
);

FILL FILL136040x232180 (
);

FILL FILL182400x345800 (
);

FILL FILL_0__14908_ (
);

FILL FILL364040x296400 (
);

OR2X2 _17665_ (
    .A(_6586_),
    .B(_6583_),
    .Y(_6587_)
);

AND2X2 _17245_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_6172_)
);

FILL FILL302480x44460 (
);

FILL FILL_0__12095_ (
);

AND2X2 _12380_ (
    .A(_2018_),
    .B(_2017_),
    .Y(_1983_[17])
);

FILL FILL_0__18741_ (
);

FILL FILL_0__18321_ (
);

FILL FILL31920x242060 (
);

DFFSR _9587_ (
    .CLK(clk_bF$buf17),
    .D(_531_[2]),
    .Q(\datapath_1.regfile_1.regOut[9] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _9167_ (
    .A(_376_),
    .B(_375_),
    .Y(_333_[21])
);

FILL FILL504640x158080 (
);

FILL FILL223440x103740 (
);

FILL FILL_0__8422_ (
);

FILL FILL_0__10408_ (
);

FILL FILL_0_BUFX2_insert870 (
);

FILL FILL_0_BUFX2_insert872 (
);

FILL FILL_0_BUFX2_insert874 (
);

INVX1 _13585_ (
    .A(PCSource[1]),
    .Y(_3080_)
);

FILL FILL_0_BUFX2_insert876 (
);

XOR2X1 _13165_ (
    .A(_2283_),
    .B(_2259_),
    .Y(_2715_)
);

FILL FILL_0_BUFX2_insert878 (
);

FILL FILL_0_BUFX2_insert879 (
);

FILL FILL_0__14661_ (
);

FILL FILL_0__14241_ (
);

FILL FILL371640x232180 (
);

FILL FILL131480x34580 (
);

FILL FILL329840x44460 (
);

FILL FILL_0__9627_ (
);

FILL FILL71440x242060 (
);

FILL FILL_1__16033_ (
);

FILL FILL_0__15866_ (
);

AND2X2 _15731_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_4682_)
);

FILL FILL_0__15026_ (
);

OR2X2 _15311_ (
    .A(_4267_),
    .B(_4266_),
    .Y(_4268_)
);

FILL FILL343520x365560 (
);

FILL FILL_0__10161_ (
);

FILL FILL326040x59280 (
);

BUFX2 BUFX2_insert30 (
    .A(_4223_),
    .Y(_4223__bF$buf4)
);

BUFX2 BUFX2_insert31 (
    .A(_4223_),
    .Y(_4223__bF$buf3)
);

BUFX2 BUFX2_insert32 (
    .A(_4223_),
    .Y(_4223__bF$buf2)
);

BUFX2 BUFX2_insert33 (
    .A(_4223_),
    .Y(_4223__bF$buf1)
);

BUFX2 BUFX2_insert34 (
    .A(_4223_),
    .Y(_4223__bF$buf0)
);

BUFX2 BUFX2_insert35 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf4 )
);

BUFX2 BUFX2_insert36 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf3 )
);

BUFX2 BUFX2_insert37 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf2 )
);

BUFX2 BUFX2_insert38 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf1 )
);

BUFX2 BUFX2_insert39 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf0 )
);

FILL FILL158840x34580 (
);

FILL FILL_1__12793_ (
);

FILL FILL_1__12373_ (
);

OR2X2 _16936_ (
    .A(_5860_),
    .B(_5867_),
    .Y(_5868_)
);

OR2X2 _16516_ (
    .A(_5452_),
    .B(_5453_),
    .Y(_5454_)
);

FILL FILL_0__11366_ (
);

DFFSR _11651_ (
    .CLK(clk_bF$buf112),
    .D(_1587_[2]),
    .Q(\datapath_1.regfile_1.regOut[25] [2]),
    .R(rst_bF$buf3),
    .S(vdd)
);

AND2X2 _11231_ (
    .A(_1432_),
    .B(_1431_),
    .Y(_1389_[21])
);

AND2X2 _8858_ (
    .A(_210_),
    .B(_209_),
    .Y(_201_[4])
);

BUFX2 _8438_ (
    .A(_2_[14]),
    .Y(memoryWriteData[14])
);

FILL FILL75240x350740 (
);

FILL FILL389880x301340 (
);

FILL FILL_1__13158_ (
);

NAND2X1 _12856_ (
    .A(_2246_),
    .B(_2420_),
    .Y(_2421_)
);

DFFSR _12436_ (
    .CLK(clk_bF$buf103),
    .D(_1983_[13]),
    .Q(\datapath_1.regfile_1.regOut[31] [13]),
    .R(rst_bF$buf32),
    .S(vdd)
);

OR2X2 _12016_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .B(_1850__bF$buf1),
    .Y(_1836_)
);

FILL FILL_0__13932_ (
);

FILL FILL_1__9121_ (
);

FILL FILL410400x44460 (
);

FILL FILL_1__15724_ (
);

FILL FILL_0__14717_ (
);

FILL FILL247760x83980 (
);

OR2X2 _17894_ (
    .A(_6804_),
    .B(_6811_),
    .Y(_6812_)
);

OR2X2 _17474_ (
    .A(_6365_),
    .B(_6398_),
    .Y(_6399_)
);

FILL FILL_0__17189_ (
);

AND2X2 _17054_ (
    .A(_4175__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_5984_)
);

FILL FILL127680x247000 (
);

FILL FILL_0__18970_ (
);

FILL FILL_0__18550_ (
);

FILL FILL350360x118560 (
);

FILL FILL_1__16929_ (
);

OR2X2 _9396_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_489_)
);

FILL FILL468160x242060 (
);

FILL FILL_1__11644_ (
);

AND2X2 _10922_ (
    .A(_1266_),
    .B(_1265_),
    .Y(_1257_[4])
);

DFFSR _10502_ (
    .CLK(clk_bF$buf47),
    .D(_993_[14]),
    .Q(\datapath_1.regfile_1.regOut[16] [14]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL35720x256880 (
);

OR2X2 _18679_ (
    .A(_7583_),
    .B(_7584_),
    .Y(_7585_)
);

AND2X2 _18259_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_7171_)
);

FILL FILL373160x202540 (
);

OAI21X1 _13394_ (
    .A(_2930_),
    .B(_2391_),
    .C(_2929_),
    .Y(_2931_)
);

FILL FILL110200x182780 (
);

FILL FILL_0__19335_ (
);

AND2X2 _19200_ (
    .A(_6232__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_8098_)
);

FILL FILL_0__14890_ (
);

FILL FILL_0__14050_ (
);

FILL FILL_0__9436_ (
);

FILL FILL_0__9016_ (
);

OR2X2 _11707_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .B(_1718__bF$buf3),
    .Y(_1670_)
);

FILL FILL284240x365560 (
);

DFFSR _14599_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[5]),
    .Q(\aluControl_1.inst [5]),
    .R(rst_bF$buf100),
    .S(vdd)
);

FILL FILL324520x79040 (
);

OR2X2 _14179_ (
    .A(MemToReg_bF$buf0),
    .B(ALUOut[12]),
    .Y(_3564_)
);

FILL FILL_1__16682_ (
);

OR2X2 _15960_ (
    .A(_4906_),
    .B(_4899_),
    .Y(_4907_)
);

FILL FILL_0__15675_ (
);

AND2X2 _15540_ (
    .A(_4142__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_4494_)
);

FILL FILL_0__15255_ (
);

NAND2X1 _15120_ (
    .A(_4017_),
    .B(_4013_),
    .Y(_4098_)
);

FILL FILL298680x326040 (
);

FILL FILL_1__17047_ (
);

OR2X2 _10099_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .B(_860__bF$buf1),
    .Y(_858_)
);

AND2X2 _16745_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_5680_)
);

AND2X2 _16325_ (
    .A(_4195__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_5266_)
);

FILL FILL_0__11595_ (
);

OR2X2 _11880_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_1765_)
);

OR2X2 _11460_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_1545_)
);

FILL FILL_0__11175_ (
);

FILL FILL436240x54340 (
);

OR2X2 _11040_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_1325_)
);

FILL FILL170240x19760 (
);

FILL FILL_0__17821_ (
);

FILL FILL12160x64220 (
);

OR2X2 _8667_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_123_)
);

FILL FILL314640x266760 (
);

INVX1 _12665_ (
    .A(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2230_)
);

AND2X2 _12245_ (
    .A(_1948_),
    .B(_1947_),
    .Y(_1917_[15])
);

FILL FILL_0__13741_ (
);

FILL FILL_0__13321_ (
);

FILL FILL195320x316160 (
);

FILL FILL282720x321100 (
);

FILL FILL39520x64220 (
);

OR2X2 _14811_ (
    .A(\datapath_1.rd2 [18]),
    .B(_3935__bF$buf4),
    .Y(_3907_)
);

FILL FILL_0__14526_ (
);

FILL FILL_0__14106_ (
);

FILL FILL354160x0 (
);

AND2X2 _17283_ (
    .A(_6208_),
    .B(\datapath_1.PCJump [26]),
    .Y(_6209_)
);

FILL FILL63840x261820 (
);

FILL FILL82080x330980 (
);

FILL FILL_1__11453_ (
);

FILL FILL367840x172900 (
);

FILL FILL_0__8880_ (
);

FILL FILL_0__10866_ (
);

FILL FILL_0__10446_ (
);

OR2X2 _10731_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_1179_)
);

OR2X2 _10311_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_959_)
);

OR2X2 _18488_ (
    .A(_7393_),
    .B(_7396_),
    .Y(_7397_)
);

OR2X2 _18068_ (
    .A(_6978_),
    .B(_6982_),
    .Y(_6983_)
);

FILL FILL297920x177840 (
);

FILL FILL_0__19144_ (
);

FILL FILL_1__12658_ (
);

FILL FILL_0__9245_ (
);

DFFSR _11936_ (
    .CLK(clk_bF$buf53),
    .D(_1719_[29]),
    .Q(\datapath_1.regfile_1.regOut[27] [29]),
    .R(rst_bF$buf111),
    .S(vdd)
);

AND2X2 _11516_ (
    .A(_1582_),
    .B(_1581_),
    .Y(_1521_[30])
);

FILL FILL132240x49400 (
);

FILL FILL_1__16071_ (
);

FILL FILL37240x88920 (
);

FILL FILL_1_BUFX2_insert90 (
);

FILL FILL_1_BUFX2_insert92 (
);

FILL FILL_1__17696_ (
);

FILL FILL_0__16689_ (
);

AND2X2 _16974_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_5905_)
);

AND2X2 _16554_ (
    .A(_4146__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_5492_)
);

FILL FILL_0__16269_ (
);

FILL FILL183160x83980 (
);

AND2X2 _16134_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_5078_)
);

FILL FILL386840x158080 (
);

FILL FILL_1__9406_ (
);

FILL FILL_0__17630_ (
);

FILL FILL_0__17210_ (
);

FILL FILL55480x182780 (
);

OR2X2 _8896_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .B(_266__bF$buf1),
    .Y(_236_)
);

OR2X2 _8476_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .B(_68__bF$buf3),
    .Y(_16_)
);

FILL FILL424080x9880 (
);

FILL FILL_1__10724_ (
);

OR2X2 _17759_ (
    .A(_6678_),
    .B(_6677_),
    .Y(_6679_)
);

AND2X2 _17339_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_6265_)
);

AOI22X1 _12894_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .C(\datapath_1.alu_1.ALUInA [16]),
    .D(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2459_)
);

INVX1 _12474_ (
    .A(\aluControl_1.inst [5]),
    .Y(_2067_)
);

DFFSR _12054_ (
    .CLK(clk_bF$buf67),
    .D(_1785_[18]),
    .Q(\datapath_1.regfile_1.regOut[28] [18]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL259160x187720 (
);

FILL FILL_0__18835_ (
);

AND2X2 _18700_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_7606_)
);

FILL FILL_0__18415_ (
);

FILL FILL_0__13550_ (
);

FILL FILL_0__13130_ (
);

FILL FILL_0__8516_ (
);

FILL FILL276640x197600 (
);

FILL FILL_1_BUFX2_insert1180 (
);

FILL FILL_1_BUFX2_insert1182 (
);

AND2X2 _13679_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3162_)
);

AND2X2 _13259_ (
    .A(_2803_),
    .B(_2800_),
    .Y(_2804_)
);

DFFSR _14620_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[26]),
    .Q(\control_1.op [0]),
    .R(rst_bF$buf100),
    .S(vdd)
);

FILL FILL425600x182780 (
);

OR2X2 _14200_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[19]),
    .Y(_3578_)
);

FILL FILL462080x9880 (
);

OR2X2 _17092_ (
    .A(_6019_),
    .B(_6020_),
    .Y(_6021_)
);

FILL FILL491720x14820 (
);

FILL FILL_1__16547_ (
);

FILL FILL432440x98800 (
);

FILL FILL503880x291460 (
);

FILL FILL414960x69160 (
);

AND2X2 _15825_ (
    .A(_4183__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_4774_)
);

AND2X2 _15405_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_4361_)
);

FILL FILL_0__10675_ (
);

OR2X2 _10960_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .B(_1322__bF$buf3),
    .Y(_1292_)
);

OR2X2 _10540_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .B(_1124__bF$buf3),
    .Y(_1072_)
);

DFFSR _10120_ (
    .CLK(clk_bF$buf60),
    .D(_795_[19]),
    .Q(\datapath_1.regfile_1.regOut[13] [19]),
    .R(rst_bF$buf59),
    .S(vdd)
);

AND2X2 _18297_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_7209_)
);

FILL FILL183920x227240 (
);

FILL FILL_1__12887_ (
);

FILL FILL_0__9894_ (
);

OR2X2 _11745_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_1695_)
);

FILL FILL_0__9054_ (
);

OR2X2 _11325_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_1475_)
);

FILL FILL261440x88920 (
);

FILL FILL_0__12821_ (
);

FILL FILL_0__15293_ (
);

FILL FILL_0__13606_ (
);

FILL FILL69160x4940 (
);

FILL FILL_0__16498_ (
);

OR2X2 _16783_ (
    .A(_5715_),
    .B(_5716_),
    .Y(_5717_)
);

FILL FILL_0__16078_ (
);

OR2X2 _16363_ (
    .A(_5303_),
    .B(_5302_),
    .Y(_5304_)
);

FILL FILL219640x202540 (
);

FILL FILL_1__10533_ (
);

BUFX2 BUFX2_insert470 (
    .A(_1388_),
    .Y(_1388__bF$buf0)
);

BUFX2 BUFX2_insert471 (
    .A(_6312_),
    .Y(_6312__bF$buf4)
);

BUFX2 BUFX2_insert472 (
    .A(_6312_),
    .Y(_6312__bF$buf3)
);

BUFX2 BUFX2_insert473 (
    .A(_6312_),
    .Y(_6312__bF$buf2)
);

BUFX2 BUFX2_insert474 (
    .A(_6312_),
    .Y(_6312__bF$buf1)
);

AND2X2 _17988_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_6905_)
);

OR2X2 _17568_ (
    .A(_6483_),
    .B(_6490_),
    .Y(_6491_)
);

BUFX2 BUFX2_insert475 (
    .A(_6312_),
    .Y(_6312__bF$buf0)
);

BUFX2 BUFX2_insert476 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf4 )
);

AND2X2 _17148_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_6076_)
);

BUFX2 BUFX2_insert477 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf3 )
);

BUFX2 BUFX2_insert478 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf2 )
);

BUFX2 BUFX2_insert479 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf1 )
);

OR2X2 _12283_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .B(_1982__bF$buf2),
    .Y(_1974_)
);

FILL FILL_1__19231_ (
);

FILL FILL_0__18644_ (
);

FILL FILL_0__8745_ (
);

OR2X2 _13488_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .B(IorD_bF$buf3),
    .Y(_3078_)
);

XOR2X1 _13068_ (
    .A(_2264_),
    .B(_2603_),
    .Y(_2624_)
);

FILL FILL_1__15151_ (
);

FILL FILL_0__19429_ (
);

FILL FILL_0__19009_ (
);

FILL FILL_0__14564_ (
);

FILL FILL_0__14144_ (
);

FILL FILL76000x330980 (
);

FILL FILL454480x108680 (
);

FILL FILL48640x365560 (
);

FILL FILL_0__15769_ (
);

FILL FILL_0__15349_ (
);

AND2X2 _15634_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_4586_)
);

AND2X2 _15214_ (
    .A(_4169_),
    .B(_4171_),
    .Y(_4172_)
);

FILL FILL_0__10484_ (
);

FILL FILL_0__10064_ (
);

FILL FILL_0__16710_ (
);

FILL FILL447640x9880 (
);

FILL FILL196840x266760 (
);

FILL FILL124640x306280 (
);

FILL FILL_0__19182_ (
);

FILL FILL11400x108680 (
);

OR2X2 _16839_ (
    .A(_5771_),
    .B(_5770_),
    .Y(_5772_)
);

OR2X2 _16419_ (
    .A(_5358_),
    .B(_5357_),
    .Y(_5359_)
);

OR2X2 _11974_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_1850__bF$buf3),
    .Y(_1808_)
);

FILL FILL_0__9283_ (
);

OR2X2 _11554_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(_1652__bF$buf0),
    .Y(_1588_)
);

DFFSR _11134_ (
    .CLK(clk_bF$buf1),
    .D(_1323_[1]),
    .Q(\datapath_1.regfile_1.regOut[21] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL_0__17915_ (
);

FILL FILL277400x133380 (
);

FILL FILL_0__12210_ (
);

FILL FILL433960x39520 (
);

FILL FILL60040x133380 (
);

FILL FILL446120x9880 (
);

OR2X2 _9702_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_653_)
);

FILL FILL97280x256880 (
);

NOR2X1 _12759_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2324_)
);

OR2X2 _12339_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_1991_)
);

FILL FILL_1__14842_ (
);

FILL FILL449920x4940 (
);

FILL FILL_0__13415_ (
);

AND2X2 _13700_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3180_)
);

FILL FILL19000x271700 (
);

OR2X2 _16592_ (
    .A(_5525_),
    .B(_5528_),
    .Y(_5529_)
);

AND2X2 _16172_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_5116_)
);

FILL FILL440040x34580 (
);

FILL FILL_1__9444_ (
);

FILL FILL_1__10342_ (
);

AND2X2 _14905_ (
    .A(_3949_),
    .B(_3948_),
    .Y(_3936_[6])
);

FILL FILL46360x227240 (
);

FILL FILL177080x118560 (
);

OR2X2 _17797_ (
    .A(_6701_),
    .B(_6716_),
    .Y(_6717_)
);

AND2X2 _17377_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_6303_)
);

FILL FILL_1__19460_ (
);

AND2X2 _12092_ (
    .A(_1866_),
    .B(_1865_),
    .Y(_1851_[7])
);

FILL FILL_0__18453_ (
);

FILL FILL_0__18033_ (
);

AND2X2 _9299_ (
    .A(_444_),
    .B(_443_),
    .Y(_399_[22])
);

FILL FILL467400x34580 (
);

FILL FILL_0__8974_ (
);

OR2X2 _10825_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .B(_1256__bF$buf4),
    .Y(_1222_)
);

OR2X2 _10405_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_1058__bF$buf1),
    .Y(_1002_)
);

NAND3X1 _13297_ (
    .A(_2383_),
    .B(ALUControl[1]),
    .C(_2425_),
    .Y(_2839_)
);

DFFSR _19523_ (
    .CLK(clk_bF$buf105),
    .D(_8320_[0]),
    .Q(\datapath_1.regfile_1.regOut[0] [0]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL_0__19238_ (
);

OR2X2 _19103_ (
    .A(_8001_),
    .B(_8000_),
    .Y(_8002_)
);

FILL FILL_0__14793_ (
);

FILL FILL_0__14373_ (
);

FILL FILL243200x207480 (
);

FILL FILL110200x296400 (
);

FILL FILL399760x123500 (
);

FILL FILL107160x247000 (
);

FILL FILL_0__9759_ (
);

FILL FILL338960x232180 (
);

FILL FILL_1__16165_ (
);

FILL FILL186200x158080 (
);

FILL FILL505400x49400 (
);

FILL FILL_0__15998_ (
);

FILL FILL247000x128440 (
);

OR2X2 _15863_ (
    .A(_4804_),
    .B(_4811_),
    .Y(_4812_)
);

FILL FILL207480x340860 (
);

FILL FILL_0__15158_ (
);

OR2X2 _15443_ (
    .A(_4396_),
    .B(_4397_),
    .Y(_4398_)
);

XOR2X1 _15023_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_4012_)
);

FILL FILL_0__10293_ (
);

FILL FILL228000x286520 (
);

FILL FILL224960x350740 (
);

FILL FILL325280x237120 (
);

OR2X2 _16648_ (
    .A(_5580_),
    .B(_5583_),
    .Y(_5584_)
);

AND2X2 _16228_ (
    .A(_4208__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_5171_)
);

FILL FILL_0__11498_ (
);

DFFSR _11783_ (
    .CLK(clk_bF$buf7),
    .D(_1653_[5]),
    .Q(\datapath_1.regfile_1.regOut[26] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL_1__18311_ (
);

AND2X2 _11363_ (
    .A(_1500_),
    .B(_1499_),
    .Y(_1455_[22])
);

FILL FILL_0__17304_ (
);

FILL FILL348080x321100 (
);

FILL FILL241680x266760 (
);

FILL FILL281200x375440 (
);

FILL FILL204440x0 (
);

OR2X2 _9931_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .B(_794__bF$buf2),
    .Y(_766_)
);

OR2X2 _9511_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .B(_596__bF$buf3),
    .Y(_546_)
);

AOI22X1 _12988_ (
    .A(_2323_),
    .B(_2379__bF$buf3),
    .C(_2548_),
    .D(_2324_),
    .Y(_2549_)
);

OR2X2 _12568_ (
    .A(_2079_),
    .B(_2088_),
    .Y(_2089_)
);

OR2X2 _12148_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .B(_1916__bF$buf1),
    .Y(_1904_)
);

FILL FILL_0__18929_ (
);

FILL FILL_0__18509_ (
);

FILL FILL104120x330980 (
);

FILL FILL107920x98800 (
);

FILL FILL_0__13644_ (
);

FILL FILL_0__13224_ (
);

FILL FILL_1__9253_ (
);

BUFX2 BUFX2_insert1030 (
    .A(_662_),
    .Y(_662__bF$buf4)
);

BUFX2 BUFX2_insert1031 (
    .A(_662_),
    .Y(_662__bF$buf3)
);

BUFX2 BUFX2_insert1032 (
    .A(_662_),
    .Y(_662__bF$buf2)
);

BUFX2 BUFX2_insert1033 (
    .A(_662_),
    .Y(_662__bF$buf1)
);

BUFX2 BUFX2_insert1034 (
    .A(_662_),
    .Y(_662__bF$buf0)
);

BUFX2 BUFX2_insert1035 (
    .A(_6272_),
    .Y(_6272__bF$buf4)
);

BUFX2 BUFX2_insert1036 (
    .A(_6272_),
    .Y(_6272__bF$buf3)
);

BUFX2 BUFX2_insert1037 (
    .A(_6272_),
    .Y(_6272__bF$buf2)
);

BUFX2 BUFX2_insert1038 (
    .A(_6272_),
    .Y(_6272__bF$buf1)
);

FILL FILL_1__15016_ (
);

BUFX2 BUFX2_insert1039 (
    .A(_6272_),
    .Y(_6272__bF$buf0)
);

FILL FILL_1__10151_ (
);

FILL FILL_0__14849_ (
);

OR2X2 _14714_ (
    .A(vdd),
    .B(\datapath_1.a [29]),
    .Y(_3862_)
);

FILL FILL_0__14429_ (
);

FILL FILL_0__14009_ (
);

BUFX2 BUFX2_insert850 (
    .A(_6317_),
    .Y(_6317__bF$buf2)
);

BUFX2 BUFX2_insert851 (
    .A(_6317_),
    .Y(_6317__bF$buf1)
);

BUFX2 BUFX2_insert852 (
    .A(_6317_),
    .Y(_6317__bF$buf0)
);

BUFX2 BUFX2_insert853 (
    .A(_4001_),
    .Y(_4001__bF$buf4)
);

BUFX2 BUFX2_insert854 (
    .A(_4001_),
    .Y(_4001__bF$buf3)
);

BUFX2 BUFX2_insert855 (
    .A(_4001_),
    .Y(_4001__bF$buf2)
);

BUFX2 BUFX2_insert856 (
    .A(_4001_),
    .Y(_4001__bF$buf1)
);

AND2X2 _17186_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_6114_)
);

BUFX2 BUFX2_insert857 (
    .A(_4001_),
    .Y(_4001__bF$buf0)
);

BUFX2 BUFX2_insert858 (
    .A(_4230_),
    .Y(_4230__bF$buf4)
);

BUFX2 BUFX2_insert859 (
    .A(_4230_),
    .Y(_4230__bF$buf3)
);

FILL FILL_0__18682_ (
);

FILL FILL161880x242060 (
);

FILL FILL_0__18262_ (
);

FILL FILL_1__11776_ (
);

FILL FILL457520x133380 (
);

OR2X2 _15919_ (
    .A(_4866_),
    .B(_4863_),
    .Y(_4867_)
);

FILL FILL116280x365560 (
);

FILL FILL_0__10349_ (
);

DFFSR _10634_ (
    .CLK(clk_bF$buf35),
    .D(_1059_[17]),
    .Q(\datapath_1.regfile_1.regOut[17] [17]),
    .R(rst_bF$buf6),
    .S(vdd)
);

FILL FILL6080x54340 (
);

AND2X2 _10214_ (
    .A(_914_),
    .B(_913_),
    .Y(_861_[26])
);

FILL FILL49400x24700 (
);

FILL FILL_0__19467_ (
);

OR2X2 _19332_ (
    .A(_8227_),
    .B(_8226_),
    .Y(_8228_)
);

FILL FILL_0__14182_ (
);

FILL FILL279680x232180 (
);

FILL FILL_0__9568_ (
);

OR2X2 _11839_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .B(_1784__bF$buf0),
    .Y(_1738_)
);

FILL FILL_0__9148_ (
);

DFFSR _11419_ (
    .CLK(clk_bF$buf74),
    .D(_1455_[28]),
    .Q(\datapath_1.regfile_1.regOut[23] [28]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL_0__12915_ (
);

FILL FILL_0__15387_ (
);

OR2X2 _15672_ (
    .A(_4623_),
    .B(_4608_),
    .Y(_4624_)
);

AND2X2 _15252_ (
    .A(_4157_),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_4210_)
);

FILL FILL26600x98800 (
);

FILL FILL60800x271700 (
);

FILL FILL51680x375440 (
);

AND2X2 _16877_ (
    .A(_4239__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_5810_)
);

OR2X2 _16457_ (
    .A(_5388_),
    .B(_5395_),
    .Y(_5396_)
);

FILL FILL301720x113620 (
);

AND2X2 _16037_ (
    .A(_4210__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_4983_)
);

FILL FILL_1__18960_ (
);

OR2X2 _11592_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_1613_)
);

OR2X2 _11172_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_1393_)
);

FILL FILL_0__17533_ (
);

FILL FILL218880x34580 (
);

OR2X2 _8799_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_191_)
);

DFFSR _9740_ (
    .CLK(clk_bF$buf86),
    .D(_597_[26]),
    .Q(\datapath_1.regfile_1.regOut[10] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

AND2X2 _9320_ (
    .A(_458_),
    .B(_457_),
    .Y(_399_[29])
);

FILL FILL_1__13099_ (
);

INVX1 _12797_ (
    .A(_2361_),
    .Y(_2362_)
);

FILL FILL_1__19325_ (
);

AND2X2 _12377_ (
    .A(_2016_),
    .B(_2015_),
    .Y(_1983_[16])
);

FILL FILL84360x24700 (
);

FILL FILL383800x93860 (
);

FILL FILL_1__14040_ (
);

FILL FILL_0__18318_ (
);

AND2X2 _18603_ (
    .A(_6317__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_7510_)
);

FILL FILL468160x64220 (
);

FILL FILL_0__13873_ (
);

FILL FILL148200x355680 (
);

FILL FILL197600x153140 (
);

FILL FILL_1__15665_ (
);

OR2X2 _14943_ (
    .A(\datapath_1.mux_pcsrc.dout [19]),
    .B(_4001__bF$buf0),
    .Y(_3975_)
);

FILL FILL_0__14658_ (
);

FILL FILL_0__14238_ (
);

OR2X2 _14523_ (
    .A(memoryOutData[8]),
    .B(_3803__bF$buf3),
    .Y(_3755_)
);

AND2X2 _14103_ (
    .A(_3350__bF$buf0),
    .B(_2_[26]),
    .Y(_3508_)
);

FILL FILL_0__18491_ (
);

FILL FILL_0__18071_ (
);

FILL FILL88160x24700 (
);

FILL FILL_1__11585_ (
);

AND2X2 _15728_ (
    .A(_4234__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_4679_)
);

OR2X2 _15308_ (
    .A(_4263_),
    .B(_4264_),
    .Y(_4265_)
);

FILL FILL_0__10998_ (
);

OR2X2 _10863_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_1247_)
);

FILL FILL_0__10578_ (
);

FILL FILL_1__17811_ (
);

FILL FILL_0__10158_ (
);

OR2X2 _10443_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_1027_)
);

OR2X2 _10023_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_807_)
);

FILL FILL_0__16804_ (
);

FILL FILL83600x365560 (
);

FILL FILL_0__19276_ (
);

AND2X2 _19141_ (
    .A(_6211__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_8040_)
);

FILL FILL298680x212420 (
);

FILL FILL315400x316160 (
);

FILL FILL402800x321100 (
);

FILL FILL_0__9377_ (
);

AND2X2 _11648_ (
    .A(_1650_),
    .B(_1649_),
    .Y(_1587_[31])
);

AND2X2 _11228_ (
    .A(_1430_),
    .B(_1429_),
    .Y(_1389_[20])
);

FILL FILL301720x340860 (
);

FILL FILL_0__12724_ (
);

OR2X2 _15481_ (
    .A(_4404_),
    .B(_4435_),
    .Y(_4436_)
);

FILL FILL_0__15196_ (
);

NAND2X1 _15061_ (
    .A(_4002_),
    .B(_4049_),
    .Y(_4050_)
);

FILL FILL8360x9880 (
);

FILL FILL401280x29640 (
);

FILL FILL_0__13509_ (
);

FILL FILL419520x330980 (
);

OR2X2 _16686_ (
    .A(_5621_),
    .B(_5620_),
    .Y(_5622_)
);

AND2X2 _16266_ (
    .A(_4228__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_5208_)
);

FILL FILL_1__9538_ (
);

FILL FILL_0__17762_ (
);

FILL FILL500840x167960 (
);

DFFSR _12186_ (
    .CLK(clk_bF$buf4),
    .D(_1851_[21]),
    .Q(\datapath_1.regfile_1.regOut[29] [21]),
    .R(rst_bF$buf20),
    .S(vdd)
);

FILL FILL300200x9880 (
);

FILL FILL_0__18967_ (
);

AND2X2 _18832_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_7736_)
);

FILL FILL_0__18127_ (
);

OR2X2 _18412_ (
    .A(_7321_),
    .B(_7318_),
    .Y(_7322_)
);

FILL FILL_0__13262_ (
);

FILL FILL293360x182780 (
);

FILL FILL_0__8648_ (
);

AND2X2 _10919_ (
    .A(_1264_),
    .B(_1263_),
    .Y(_1257_[3])
);

FILL FILL366320x296400 (
);

DFFSR _14752_ (
    .CLK(clk_bF$buf15),
    .D(_3804_[29]),
    .Q(\datapath_1.a [29]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL_0__14047_ (
);

AND2X2 _14332_ (
    .A(_3667_),
    .B(_3666_),
    .Y(_3606_[30])
);

FILL FILL415720x83980 (
);

FILL FILL225720x103740 (
);

AND2X2 _15957_ (
    .A(_4146__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_4904_)
);

AND2X2 _15537_ (
    .A(_4130__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_4491_)
);

AND2X2 _15117_ (
    .A(_4036_),
    .B(_4091_),
    .Y(_4096_)
);

FILL FILL142120x247000 (
);

OR2X2 _10672_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .B(_1190__bF$buf4),
    .Y(_1140_)
);

DFFSR _10252_ (
    .CLK(clk_bF$buf25),
    .D(_861_[22]),
    .Q(\datapath_1.regfile_1.regOut[14] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

FILL FILL_0__16613_ (
);

FILL FILL373920x232180 (
);

OR2X2 _19370_ (
    .A(_8264_),
    .B(_8263_),
    .Y(_8265_)
);

DFFSR _8820_ (
    .CLK(clk_bF$buf102),
    .D(_135_[9]),
    .Q(\datapath_1.regfile_1.regOut[3] [9]),
    .R(rst_bF$buf59),
    .S(vdd)
);

BUFX2 _8400_ (
    .A(_1_[8]),
    .Y(memoryAddress[8])
);

FILL FILL424080x291460 (
);

FILL FILL415720x360620 (
);

FILL FILL73720x242060 (
);

FILL FILL305520x14820 (
);

FILL FILL159600x350740 (
);

FILL FILL_1__18825_ (
);

OR2X2 _11877_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_1763_)
);

FILL FILL_0__9186_ (
);

OR2X2 _11457_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_1543_)
);

INVX2 _11037_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .Y(_1388_)
);

FILL FILL_1__13540_ (
);

FILL FILL256880x301340 (
);

FILL FILL_0__12533_ (
);

FILL FILL345800x365560 (
);

FILL FILL_0__12113_ (
);

FILL FILL215840x49400 (
);

AND2X2 _15290_ (
    .A(_4247_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd2 [0])
);

DFFSR _9605_ (
    .CLK(clk_bF$buf9),
    .D(_531_[20]),
    .Q(\datapath_1.regfile_1.regOut[9] [20]),
    .R(rst_bF$buf28),
    .S(vdd)
);

FILL FILL383040x321100 (
);

FILL FILL_0__13738_ (
);

OR2X2 _13603_ (
    .A(_3096_),
    .B(_3095_),
    .Y(_3097_)
);

OR2X2 _16495_ (
    .A(_5430_),
    .B(_5433_),
    .Y(_5434_)
);

AND2X2 _16075_ (
    .A(_4167__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_5020_)
);

FILL FILL_0__17571_ (
);

FILL FILL112480x64220 (
);

FILL FILL_0__17151_ (
);

FILL FILL77520x350740 (
);

FILL FILL464360x251940 (
);

OR2X2 _14808_ (
    .A(\datapath_1.rd2 [17]),
    .B(_3935__bF$buf0),
    .Y(_3905_)
);

FILL FILL309320x301340 (
);

FILL FILL96520x34580 (
);

FILL FILL_0__18776_ (
);

OR2X2 _18641_ (
    .A(_7540_),
    .B(_7547_),
    .Y(_7548_)
);

FILL FILL_0__18356_ (
);

AND2X2 _18221_ (
    .A(_6259__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_7134_)
);

FILL FILL_0__13491_ (
);

FILL FILL_0__8877_ (
);

FILL FILL_0__8457_ (
);

OR2X2 _10728_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_1177_)
);

FILL FILL433200x44460 (
);

OR2X2 _10308_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_957_)
);

FILL FILL_1__15283_ (
);

OR2X2 _19426_ (
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .B(gnd),
    .Y(_8384_)
);

OR2X2 _19006_ (
    .A(_7905_),
    .B(_7906_),
    .Y(_7907_)
);

FILL FILL138320x370500 (
);

DFFSR _14981_ (
    .CLK(clk_bF$buf62),
    .D(_3936_[0]),
    .Q(\datapath_1.mux_iord.din0 [0]),
    .R(rst_bF$buf18),
    .S(vdd)
);

FILL FILL343520x79040 (
);

OR2X2 _14561_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump [23]),
    .Y(_3780_)
);

OR2X2 _14141_ (
    .A(_3540_),
    .B(_3537_),
    .Y(\datapath_1.alu_1.ALUInB [31])
);

FILL FILL129960x247000 (
);

FILL FILL352640x118560 (
);

FILL FILL_1__16488_ (
);

OR2X2 _15766_ (
    .A(_4714_),
    .B(_4715_),
    .Y(_4716_)
);

OR2X2 _15346_ (
    .A(_4301_),
    .B(_4302_),
    .Y(_4303_)
);

FILL FILL155040x286520 (
);

FILL FILL_0__10196_ (
);

AND2X2 _10481_ (
    .A(_1052_),
    .B(_1051_),
    .Y(_993_[29])
);

AND2X2 _10061_ (
    .A(_832_),
    .B(_831_),
    .Y(_795_[18])
);

FILL FILL_0__16002_ (
);

FILL FILL47880x247000 (
);

OR2X2 _11686_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .B(_1718__bF$buf1),
    .Y(_1656_)
);

DFFSR _11266_ (
    .CLK(clk_bF$buf79),
    .D(_1389_[4]),
    .Q(\datapath_1.regfile_1.regOut[22] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL_0__17627_ (
);

AND2X2 _17912_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_6830_)
);

FILL FILL_0__12762_ (
);

FILL FILL_0__12342_ (
);

FILL FILL132240x311220 (
);

OR2X2 _9834_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_721_)
);

OR2X2 _9414_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_501_)
);

FILL FILL_1__14974_ (
);

FILL FILL_0__13967_ (
);

OR2X2 _13832_ (
    .A(\datapath_1.a [5]),
    .B(_3342__bF$buf2),
    .Y(_3288_)
);

FILL FILL_0__13127_ (
);

AND2X2 _13412_ (
    .A(_2945_),
    .B(_2947_),
    .Y(_2948_)
);

FILL FILL459040x54340 (
);

FILL FILL90440x296400 (
);

FILL FILL230280x291460 (
);

FILL FILL_1__9156_ (
);

FILL FILL_0__17380_ (
);

FILL FILL_1__10474_ (
);

DFFSR _14617_ (
    .CLK(clk_bF$buf11),
    .D(_3738_[23]),
    .Q(\datapath_1.PCJump [25]),
    .R(rst_bF$buf26),
    .S(vdd)
);

FILL FILL495520x44460 (
);

OR2X2 _17089_ (
    .A(_6014_),
    .B(_6017_),
    .Y(_6018_)
);

FILL FILL197600x316160 (
);

FILL FILL16720x276640 (
);

AND2X2 _18870_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_7773_)
);

FILL FILL_0__18585_ (
);

AND2X2 _18450_ (
    .A(_7359_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd1 [16])
);

AND2X2 _18030_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_6946_)
);

FILL FILL234840x172900 (
);

FILL FILL284240x227240 (
);

FILL FILL_1__17905_ (
);

OR2X2 _10957_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_1322__bF$buf3),
    .Y(_1290_)
);

OR2X2 _10537_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .B(_1124__bF$buf3),
    .Y(_1070_)
);

DFFSR _10117_ (
    .CLK(clk_bF$buf5),
    .D(_795_[16]),
    .Q(\datapath_1.regfile_1.regOut[13] [16]),
    .R(rst_bF$buf112),
    .S(vdd)
);

FILL FILL494000x103740 (
);

FILL FILL_0__11613_ (
);

AND2X2 _19235_ (
    .A(_6206__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_8132_)
);

OR2X2 _14790_ (
    .A(\datapath_1.rd2 [11]),
    .B(_3935__bF$buf4),
    .Y(_3893_)
);

FILL FILL_0__14085_ (
);

OR2X2 _14370_ (
    .A(memoryOutData[0]),
    .B(_3737__bF$buf3),
    .Y(_3673_)
);

FILL FILL98040x306280 (
);

FILL FILL_1__13405_ (
);

AND2X2 _15995_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_4941_)
);

OR2X2 _15575_ (
    .A(_4524_),
    .B(_4527_),
    .Y(_4528_)
);

NAND2X1 _15155_ (
    .A(_4059_),
    .B(_4013_),
    .Y(_4119_)
);

FILL FILL300200x167960 (
);

OR2X2 _10290_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_945_)
);

FILL FILL_1__8847_ (
);

FILL FILL_0__16651_ (
);

FILL FILL_0__16231_ (
);

FILL FILL128440x113620 (
);

FILL FILL262200x281580 (
);

AND2X2 _11495_ (
    .A(_1568_),
    .B(_1567_),
    .Y(_1521_[23])
);

AND2X2 _11075_ (
    .A(_1348_),
    .B(_1347_),
    .Y(_1323_[12])
);

FILL FILL_0__17856_ (
);

FILL FILL_0__17436_ (
);

AND2X2 _17721_ (
    .A(_6297__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_6642_)
);

NOR2X1 _17301_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_6227_)
);

FILL FILL_0__17016_ (
);

FILL FILL_0__12991_ (
);

FILL FILL_0__12571_ (
);

FILL FILL401280x360620 (
);

FILL FILL411920x59280 (
);

OR2X2 _9643_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .B(_662__bF$buf3),
    .Y(_614_)
);

DFFSR _9223_ (
    .CLK(clk_bF$buf80),
    .D(_333_[25]),
    .Q(\datapath_1.regfile_1.regOut[6] [25]),
    .R(rst_bF$buf76),
    .S(vdd)
);

FILL FILL474240x24700 (
);

FILL FILL204440x59280 (
);

AND2X2 _18926_ (
    .A(_6312__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_7828_)
);

OR2X2 _18506_ (
    .A(_7413_),
    .B(_7414_),
    .Y(_7415_)
);

FILL FILL_0__13776_ (
);

FILL FILL_0__13356_ (
);

AND2X2 _13641_ (
    .A(_3084__bF$buf4),
    .B(\aluControl_1.inst [5]),
    .Y(_3129_)
);

MUX2X1 _13221_ (
    .A(_2376__bF$buf0),
    .B(_2501_),
    .S(_2441_),
    .Y(_2768_)
);

FILL FILL57760x182780 (
);

FILL FILL_1__10283_ (
);

OR2X2 _14846_ (
    .A(vdd),
    .B(_2_[30]),
    .Y(_3930_)
);

OR2X2 _14426_ (
    .A(vdd),
    .B(\datapath_1.Data [19]),
    .Y(_3710_)
);

AND2X2 _14006_ (
    .A(_3352__bF$buf0),
    .B(\datapath_1.PCJump [12]),
    .Y(_3425_)
);

FILL FILL286520x64220 (
);

FILL FILL_0__15922_ (
);

FILL FILL_0__15502_ (
);

FILL FILL361760x187720 (
);

FILL FILL_1__11488_ (
);

FILL FILL365560x0 (
);

FILL FILL297160x266760 (
);

FILL FILL61560x197600 (
);

DFFSR _10766_ (
    .CLK(clk_bF$buf27),
    .D(_1125_[20]),
    .Q(\datapath_1.regfile_1.regOut[18] [20]),
    .R(rst_bF$buf28),
    .S(vdd)
);

AND2X2 _10346_ (
    .A(_982_),
    .B(_981_),
    .Y(_927_[27])
);

FILL FILL_0__11002_ (
);

OR2X2 _19464_ (
    .A(gnd),
    .B(_8385__bF$buf2),
    .Y(_8345_)
);

AND2X2 _19044_ (
    .A(_6272__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_7944_)
);

OR2X2 _8914_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .B(_266__bF$buf4),
    .Y(_248_)
);

FILL FILL433200x350740 (
);

FILL FILL455240x98800 (
);

FILL FILL_1__13634_ (
);

FILL FILL_1_BUFX2_insert421 (
);

INVX1 _12912_ (
    .A(_2335_),
    .Y(_2477_)
);

FILL FILL_0__12627_ (
);

FILL FILL_1_BUFX2_insert423 (
);

FILL FILL32680x281580 (
);

OR2X2 _15384_ (
    .A(_4332_),
    .B(_4339_),
    .Y(_4340_)
);

FILL FILL_0__16880_ (
);

FILL FILL_0__16040_ (
);

FILL FILL346560x330980 (
);

AND2X2 _16589_ (
    .A(_4160__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_5526_)
);

AND2X2 _16169_ (
    .A(_4177__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_5113_)
);

FILL FILL_1__18252_ (
);

FILL FILL266760x59280 (
);

OR2X2 _17950_ (
    .A(_6863_),
    .B(_6866_),
    .Y(_6867_)
);

FILL FILL_0__17245_ (
);

AND2X2 _17530_ (
    .A(_6300__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_6454_)
);

OR2X2 _17110_ (
    .A(_6037_),
    .B(_6038_),
    .Y(_6039_)
);

FILL FILL_0__12380_ (
);

FILL FILL202920x79040 (
);

FILL FILL458280x19760 (
);

DFFSR _9872_ (
    .CLK(clk_bF$buf88),
    .D(_663_[29]),
    .Q(\datapath_1.regfile_1.regOut[11] [29]),
    .R(rst_bF$buf95),
    .S(vdd)
);

AND2X2 _9452_ (
    .A(_526_),
    .B(_525_),
    .Y(_465_[30])
);

AND2X2 _9032_ (
    .A(_306_),
    .B(_305_),
    .Y(_267_[19])
);

AND2X2 _12089_ (
    .A(_1864_),
    .B(_1863_),
    .Y(_1851_[6])
);

FILL FILL_1__14592_ (
);

AND2X2 _18735_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_7640_)
);

OR2X2 _18315_ (
    .A(_7223_),
    .B(_7226_),
    .Y(_7227_)
);

OR2X2 _13870_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [18]),
    .Y(_3313_)
);

FILL FILL_0__13585_ (
);

FILL FILL_0__13165_ (
);

AND2X2 _13450_ (
    .A(_2538_),
    .B(_2571_),
    .Y(_2983_)
);

XOR2X1 _13030_ (
    .A(_2335_),
    .B(_2317_),
    .Y(_2588_)
);

FILL FILL293360x296400 (
);

FILL FILL247760x143260 (
);

OR2X2 _14655_ (
    .A(\datapath_1.rd1 [9]),
    .B(_3869__bF$buf4),
    .Y(_3823_)
);

AND2X2 _14235_ (
    .A(_3601_),
    .B(_3600_),
    .Y(\datapath_1.mux_wd3.dout [30])
);

FILL FILL107160x54340 (
);

FILL FILL_0__15731_ (
);

FILL FILL21280x83980 (
);

FILL FILL253080x311220 (
);

FILL FILL_1__17943_ (
);

OR2X2 _10995_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_1315_)
);

OR2X2 _10575_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_1095_)
);

OR2X2 _10155_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_875_)
);

FILL FILL_0__16516_ (
);

AND2X2 _16801_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_5735_)
);

AND2X2 _19273_ (
    .A(_6211__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_8170_)
);

FILL FILL318440x54340 (
);

FILL FILL190000x286520 (
);

AND2X2 _8723_ (
    .A(_140_),
    .B(_139_),
    .Y(_135_[2])
);

FILL FILL_1__13023_ (
);

FILL FILL_0__12856_ (
);

OR2X2 _12721_ (
    .A(_2276_),
    .B(_2285_),
    .Y(_2286_)
);

FILL FILL4560x247000 (
);

FILL FILL_0__12016_ (
);

DFFSR _12301_ (
    .CLK(clk_bF$buf68),
    .D(_1917_[7]),
    .Q(\datapath_1.regfile_1.regOut[30] [7]),
    .R(rst_bF$buf21),
    .S(vdd)
);

FILL FILL281960x256880 (
);

NOR3X1 _15193_ (
    .A(_4145_),
    .B(\datapath_1.PCJump_22_bF$buf0 ),
    .C(_4150_),
    .Y(_4151_)
);

OR2X2 _9928_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .B(_794__bF$buf3),
    .Y(_764_)
);

OR2X2 _9508_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .B(_596__bF$buf3),
    .Y(_544_)
);

FILL FILL126920x306280 (
);

FILL FILL323000x321100 (
);

FILL FILL_1__14648_ (
);

AND2X2 _13926_ (
    .A(_3347__bF$buf2),
    .B(\aluControl_1.inst [1]),
    .Y(_3356_)
);

AND2X2 _13506_ (
    .A(_3025_),
    .B(_3024_),
    .Y(_1_[5])
);

FILL FILL213560x217360 (
);

FILL FILL300960x222300 (
);

AND2X2 _16398_ (
    .A(_4177__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_5338_)
);

FILL FILL_0__17894_ (
);

FILL FILL_0__17474_ (
);

FILL FILL_0__17054_ (
);

FILL FILL99560x256880 (
);

OR2X2 _9681_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_639_)
);

OR2X2 _9261_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_419_)
);

FILL FILL_1_CLKBUF1_insert137 (
);

FILL FILL_1__19266_ (
);

FILL FILL_1_CLKBUF1_insert139 (
);

OR2X2 _18964_ (
    .A(_7864_),
    .B(_7865_),
    .Y(_7866_)
);

FILL FILL62320x44460 (
);

OR2X2 _18544_ (
    .A(_7444_),
    .B(_7451_),
    .Y(_7452_)
);

OR2X2 _18124_ (
    .A(_7005_),
    .B(_7038_),
    .Y(_7039_)
);

FILL FILL_0__19200_ (
);

FILL FILL374680x158080 (
);

FILL FILL_0__11707_ (
);

FILL FILL179360x118560 (
);

OR2X2 _19329_ (
    .A(_8223_),
    .B(_8224_),
    .Y(_8225_)
);

OR2X2 _14884_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .B(PCEn_bF$buf4),
    .Y(_4000_)
);

FILL FILL_0__14179_ (
);

AND2X2 _14464_ (
    .A(_3735_),
    .B(_3734_),
    .Y(_3672_[31])
);

AND2X2 _14044_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3457_)
);

FILL FILL_0__15120_ (
);

FILL FILL66120x44460 (
);

OR2X2 _15669_ (
    .A(_4620_),
    .B(_4619_),
    .Y(_4621_)
);

AND2X2 _15249_ (
    .A(_4127_),
    .B(_4139_),
    .Y(_4207_)
);

FILL FILL283480x360620 (
);

DFFSR _10384_ (
    .CLK(clk_bF$buf81),
    .D(_927_[25]),
    .Q(\datapath_1.regfile_1.regOut[15] [25]),
    .R(rst_bF$buf101),
    .S(vdd)
);

FILL FILL149720x24700 (
);

FILL FILL397480x108680 (
);

FILL FILL_0__16745_ (
);

AND2X2 _16610_ (
    .A(_4177__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_5547_)
);

FILL FILL_0__16325_ (
);

FILL FILL_0__11880_ (
);

FILL FILL_0__11460_ (
);

FILL FILL_0__11040_ (
);

FILL FILL402040x113620 (
);

AND2X2 _19082_ (
    .A(_6271__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .Y(_7982_)
);

DFFSR _8952_ (
    .CLK(clk_bF$buf113),
    .D(_201_[12]),
    .Q(\datapath_1.regfile_1.regOut[4] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

OR2X2 _8532_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_53_)
);

OR2X2 _11589_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_1611_)
);

FILL FILL_1__18117_ (
);

OR2X2 _11169_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_1391_)
);

FILL FILL78280x276640 (
);

FILL FILL323760x316160 (
);

OR2X2 _17815_ (
    .A(_6730_),
    .B(_6733_),
    .Y(_6734_)
);

FILL FILL_1_BUFX2_insert801 (
);

AND2X2 _12950_ (
    .A(_2512_),
    .B(_2357_),
    .Y(_2513_)
);

FILL FILL_1_BUFX2_insert803 (
);

FILL FILL_0__12245_ (
);

AND2X2 _12530_ (
    .A(_2119_),
    .B(\control_1.op [5]),
    .Y(_2120_)
);

AND2X2 _12110_ (
    .A(_1878_),
    .B(_1877_),
    .Y(_1851_[13])
);

DFFSR _9737_ (
    .CLK(clk_bF$buf87),
    .D(_597_[23]),
    .Q(\datapath_1.regfile_1.regOut[10] [23]),
    .R(rst_bF$buf2),
    .S(vdd)
);

AND2X2 _9317_ (
    .A(_456_),
    .B(_455_),
    .Y(_399_[28])
);

FILL FILL327560x237120 (
);

AND2X2 _13735_ (
    .A(_3089__bF$buf0),
    .B(gnd),
    .Y(_3210_)
);

FILL FILL226480x256880 (
);

OR2X2 _13315_ (
    .A(_2851_),
    .B(_2855_),
    .Y(_2856_)
);

FILL FILL353400x370500 (
);

FILL FILL381520x103740 (
);

FILL FILL_0__14811_ (
);

FILL FILL158080x138320 (
);

FILL FILL_1__9899_ (
);

FILL FILL139080x296400 (
);

OR2X2 _9490_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(_596__bF$buf4),
    .Y(_532_)
);

DFFSR _9070_ (
    .CLK(clk_bF$buf69),
    .D(_267_[1]),
    .Q(\datapath_1.regfile_1.regOut[5] [1]),
    .R(rst_bF$buf13),
    .S(vdd)
);

FILL FILL89680x133380 (
);

FILL FILL461320x54340 (
);

FILL FILL_0__10311_ (
);

OR2X2 _18773_ (
    .A(_7646_),
    .B(_7677_),
    .Y(_7678_)
);

FILL FILL_0__18488_ (
);

FILL FILL_0__18068_ (
);

AND2X2 _18353_ (
    .A(_6287__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_7264_)
);

FILL FILL296400x187720 (
);

FILL FILL_0__8589_ (
);

FILL FILL_1__12103_ (
);

FILL FILL_0__9950_ (
);

FILL FILL_0__9530_ (
);

DFFSR _11801_ (
    .CLK(clk_bF$buf101),
    .D(_1653_[23]),
    .Q(\datapath_1.regfile_1.regOut[26] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL_0__11516_ (
);

OR2X2 _19558_ (
    .A(PCWrite),
    .B(_8388_),
    .Y(_8389_)
);

FILL FILL484880x340860 (
);

AND2X2 _19138_ (
    .A(_6302__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_8037_)
);

OR2X2 _14693_ (
    .A(vdd),
    .B(\datapath_1.a [22]),
    .Y(_3848_)
);

OR2X2 _14273_ (
    .A(vdd),
    .B(ALUOut[11]),
    .Y(_3628_)
);

FILL FILL118560x365560 (
);

FILL FILL22040x98800 (
);

FILL FILL317680x19760 (
);

AND2X2 _15898_ (
    .A(_4228__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_4846_)
);

OR2X2 _15478_ (
    .A(_4432_),
    .B(_4429_),
    .Y(_4433_)
);

OR2X2 _15058_ (
    .A(_4043_),
    .B(_4046_),
    .Y(_4047_)
);

AND2X2 _10193_ (
    .A(_900_),
    .B(_899_),
    .Y(_861_[19])
);

FILL FILL_0__16974_ (
);

FILL FILL_0__16554_ (
);

FILL FILL446120x138320 (
);

OR2X2 _8761_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .B(_200__bF$buf1),
    .Y(_166_)
);

FILL FILL222680x286520 (
);

FILL FILL_1__18766_ (
);

FILL FILL_1__18346_ (
);

DFFSR _11398_ (
    .CLK(clk_bF$buf18),
    .D(_1455_[7]),
    .Q(\datapath_1.regfile_1.regOut[23] [7]),
    .R(rst_bF$buf107),
    .S(vdd)
);

FILL FILL329080x4940 (
);

AND2X2 _17624_ (
    .A(_6238__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_6546_)
);

FILL FILL_0__17339_ (
);

AND2X2 _17204_ (
    .A(_4160__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_6132_)
);

FILL FILL349600x172900 (
);

FILL FILL_0__12894_ (
);

FILL FILL_0__12474_ (
);

FILL FILL36480x365560 (
);

OR2X2 _9966_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_789_)
);

OR2X2 _9546_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_569_)
);

OR2X2 _9126_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_349_)
);

FILL FILL_0__8801_ (
);

FILL FILL348080x4940 (
);

AND2X2 _18829_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_7733_)
);

FILL FILL_0_BUFX2_insert460 (
);

FILL FILL53960x375440 (
);

AND2X2 _18409_ (
    .A(_6238__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_7319_)
);

FILL FILL_0_BUFX2_insert462 (
);

FILL FILL_0_BUFX2_insert463 (
);

AND2X2 _13964_ (
    .A(_3352__bF$buf1),
    .B(\aluControl_1.inst [4]),
    .Y(_3389_)
);

FILL FILL_0_BUFX2_insert464 (
);

FILL FILL_0__13679_ (
);

OR2X2 _13544_ (
    .A(ALUOut[18]),
    .B(_3079__bF$buf4),
    .Y(_3051_)
);

FILL FILL_0_BUFX2_insert465 (
);

INVX1 _13124_ (
    .A(_2453_),
    .Y(_2677_)
);

FILL FILL_0_BUFX2_insert466 (
);

FILL FILL_0_BUFX2_insert468 (
);

FILL FILL285000x345800 (
);

FILL FILL_1__9288_ (
);

FILL FILL_0__17092_ (
);

FILL FILL497800x167960 (
);

FILL FILL421800x19760 (
);

DFFSR _14749_ (
    .CLK(clk_bF$buf80),
    .D(_3804_[26]),
    .Q(\datapath_1.a [26]),
    .R(rst_bF$buf104),
    .S(vdd)
);

AND2X2 _14329_ (
    .A(_3665_),
    .B(_3664_),
    .Y(_3606_[29])
);

FILL FILL_1__16412_ (
);

FILL FILL301720x187720 (
);

FILL FILL104880x39520 (
);

FILL FILL_0__18297_ (
);

AND2X2 _18582_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_7489_)
);

OR2X2 _18162_ (
    .A(_7075_),
    .B(_7072_),
    .Y(_7076_)
);

FILL FILL250800x355680 (
);

FILL FILL20520x360620 (
);

FILL FILL17480x311220 (
);

FILL FILL237120x266760 (
);

FILL FILL_0__8398_ (
);

OR2X2 _10669_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .B(_1190__bF$buf4),
    .Y(_1138_)
);

DFFSR _10249_ (
    .CLK(clk_bF$buf99),
    .D(_861_[19]),
    .Q(\datapath_1.regfile_1.regOut[14] [19]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL_1__12752_ (
);

FILL FILL_0__11745_ (
);

OR2X2 _11610_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_1625_)
);

FILL FILL_0__11325_ (
);

OR2X2 _19367_ (
    .A(_8261_),
    .B(_8258_),
    .Y(_8262_)
);

FILL FILL84360x98800 (
);

AND2X2 _14082_ (
    .A(_3350__bF$buf4),
    .B(_2_[23]),
    .Y(_3490_)
);

FILL FILL360240x350740 (
);

DFFSR _8817_ (
    .CLK(clk_bF$buf59),
    .D(_135_[6]),
    .Q(\datapath_1.regfile_1.regOut[3] [6]),
    .R(rst_bF$buf92),
    .S(vdd)
);

NAND2X1 _12815_ (
    .A(_2379__bF$buf3),
    .B(_2377_),
    .Y(_2380_)
);

FILL FILL137560x345800 (
);

OR2X2 _15287_ (
    .A(_4244_),
    .B(_4233_),
    .Y(_4245_)
);

FILL FILL_1__17370_ (
);

FILL FILL_1__8979_ (
);

FILL FILL_0__16363_ (
);

FILL FILL459040x177840 (
);

AND2X2 _8990_ (
    .A(_278_),
    .B(_277_),
    .Y(_267_[5])
);

DFFSR _8570_ (
    .CLK(clk_bF$buf64),
    .D(_3_[17]),
    .Q(\datapath_1.regfile_1.regOut[1] [17]),
    .R(rst_bF$buf6),
    .S(vdd)
);

FILL FILL495520x350740 (
);

FILL FILL390640x172900 (
);

FILL FILL_1__18995_ (
);

FILL FILL500080x163020 (
);

FILL FILL355680x335920 (
);

FILL FILL_0__17988_ (
);

FILL FILL_0__17568_ (
);

OR2X2 _17853_ (
    .A(_6768_),
    .B(_6771_),
    .Y(_6772_)
);

FILL FILL148200x217360 (
);

AND2X2 _17433_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_6358_)
);

OR2X2 _17013_ (
    .A(_5942_),
    .B(_5943_),
    .Y(_5944_)
);

FILL FILL174040x158080 (
);

OR2X2 _9775_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_728__bF$buf0),
    .Y(_682_)
);

DFFSR _9355_ (
    .CLK(clk_bF$buf72),
    .D(_399_[28]),
    .Q(\datapath_1.regfile_1.regOut[7] [28]),
    .R(rst_bF$buf32),
    .S(vdd)
);

FILL FILL226480x326040 (
);

FILL FILL_1__14075_ (
);

AND2X2 _18638_ (
    .A(_6211__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_7545_)
);

OR2X2 _18218_ (
    .A(_7123_),
    .B(_7130_),
    .Y(_7131_)
);

AND2X2 _13773_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[26]),
    .Y(_3242_)
);

FILL FILL_0__13068_ (
);

OR2X2 _13353_ (
    .A(_2157__bF$buf0),
    .B(_2891_),
    .Y(_2892_)
);

FILL FILL_0__9815_ (
);

FILL FILL369360x9880 (
);

OR2X2 _14978_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.PCJump [31]),
    .Y(_3998_)
);

OR2X2 _14558_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_3778_)
);

AND2X2 _14138_ (
    .A(_3350__bF$buf4),
    .B(_2_[31]),
    .Y(_3538_)
);

FILL FILL284240x113620 (
);

FILL FILL_0__15634_ (
);

FILL FILL_0__15214_ (
);

FILL FILL295640x182780 (
);

OR2X2 _18391_ (
    .A(_7300_),
    .B(_7299_),
    .Y(_7301_)
);

FILL FILL408880x88920 (
);

FILL FILL57000x34580 (
);

DFFSR _10898_ (
    .CLK(clk_bF$buf26),
    .D(_1191_[23]),
    .Q(\datapath_1.regfile_1.regOut[19] [23]),
    .R(rst_bF$buf94),
    .S(vdd)
);

AND2X2 _10478_ (
    .A(_1050_),
    .B(_1049_),
    .Y(_993_[28])
);

AND2X2 _10058_ (
    .A(_830_),
    .B(_829_),
    .Y(_795_[17])
);

FILL FILL368600x296400 (
);

FILL FILL_0__16839_ (
);

OR2X2 _16704_ (
    .A(_5638_),
    .B(_5637_),
    .Y(_5639_)
);

FILL FILL_0__16419_ (
);

FILL FILL47880x360620 (
);

FILL FILL_0__11554_ (
);

AND2X2 _19176_ (
    .A(_6221__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_8074_)
);

FILL FILL117040x14820 (
);

OR2X2 _8626_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .B(_134__bF$buf1),
    .Y(_96_)
);

OR2X2 _17909_ (
    .A(_6826_),
    .B(_6825_),
    .Y(_6827_)
);

FILL FILL_0__12759_ (
);

XNOR2X1 _12624_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2189_)
);

FILL FILL144400x247000 (
);

FILL FILL211280x49400 (
);

OR2X2 _12204_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .Y(_1921_)
);

AND2X2 _15096_ (
    .A(_4059_),
    .B(_4020_),
    .Y(_4079_)
);

FILL FILL_0__16592_ (
);

FILL FILL_0__16172_ (
);

OR2X2 _13829_ (
    .A(\datapath_1.a [4]),
    .B(_3342__bF$buf1),
    .Y(_3286_)
);

AND2X2 _13409_ (
    .A(_2941_),
    .B(_2944_),
    .Y(_2945_)
);

FILL FILL_1__15912_ (
);

FILL FILL427880x306280 (
);

FILL FILL_0__14905_ (
);

FILL FILL_1__18384_ (
);

FILL FILL187720x291460 (
);

FILL FILL504640x271700 (
);

AND2X2 _17662_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_6584_)
);

AND2X2 _17242_ (
    .A(_4239__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_6169_)
);

FILL FILL422560x49400 (
);

AND2X2 _9584_ (
    .A(_594_),
    .B(_593_),
    .Y(_531_[31])
);

AND2X2 _9164_ (
    .A(_374_),
    .B(_373_),
    .Y(_333_[20])
);

FILL FILL_0__10825_ (
);

FILL FILL_0__10405_ (
);

OR2X2 _18867_ (
    .A(_7769_),
    .B(_7766_),
    .Y(_7770_)
);

FILL FILL_0_BUFX2_insert841 (
);

OR2X2 _18447_ (
    .A(_7341_),
    .B(_7356_),
    .Y(_7357_)
);

FILL FILL_0_BUFX2_insert842 (
);

AND2X2 _18027_ (
    .A(_6271__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_6943_)
);

FILL FILL_0_BUFX2_insert843 (
);

FILL FILL_0_BUFX2_insert844 (
);

FILL FILL_0__13297_ (
);

FILL FILL_0_BUFX2_insert845 (
);

OR2X2 _13582_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.PCJump [31]),
    .Y(_3076_)
);

AND2X2 _13162_ (
    .A(_2712_),
    .B(_2706_),
    .Y(_2713_)
);

FILL FILL_0_BUFX2_insert846 (
);

FILL FILL_0_BUFX2_insert848 (
);

FILL FILL_0__19103_ (
);

FILL FILL79800x350740 (
);

FILL FILL19000x64220 (
);

FILL FILL_1__12617_ (
);

FILL FILL_0__9624_ (
);

FILL FILL_1__15089_ (
);

OR2X2 _14787_ (
    .A(\datapath_1.rd2 [10]),
    .B(_3935__bF$buf0),
    .Y(_3891_)
);

DFFSR _14367_ (
    .CLK(clk_bF$buf50),
    .D(_3606_[31]),
    .Q(ALUOut[31]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL_0__15863_ (
);

FILL FILL_0__15443_ (
);

FILL FILL_0__15023_ (
);

FILL FILL76760x93860 (
);

OR2X2 _10287_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_943_)
);

FILL FILL_1__17235_ (
);

AND2X2 _16933_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_5865_)
);

OR2X2 _16513_ (
    .A(_5447_),
    .B(_5450_),
    .Y(_5451_)
);

FILL FILL477280x83980 (
);

FILL FILL366320x79040 (
);

FILL FILL240920x370500 (
);

FILL FILL310080x271700 (
);

AND2X2 _8855_ (
    .A(_208_),
    .B(_207_),
    .Y(_201_[3])
);

BUFX2 _8435_ (
    .A(_2_[11]),
    .Y(memoryWriteData[11])
);

FILL FILL_1__13575_ (
);

FILL FILL386080x133380 (
);

AND2X2 _17718_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_6639_)
);

XOR2X1 _12853_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2418_)
);

FILL FILL_0__12568_ (
);

FILL FILL_0__12148_ (
);

DFFSR _12433_ (
    .CLK(clk_bF$buf33),
    .D(_1983_[10]),
    .Q(\datapath_1.regfile_1.regOut[31] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

OR2X2 _12013_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .B(_1850__bF$buf0),
    .Y(_1834_)
);

OR2X2 _13638_ (
    .A(_3126_),
    .B(_3125_),
    .Y(_3127_)
);

OAI21X1 _13218_ (
    .A(_2215_),
    .B(_2744_),
    .C(_2764_),
    .Y(_2765_)
);

FILL FILL_0__14714_ (
);

FILL FILL375440x276640 (
);

FILL FILL323000x49400 (
);

AND2X2 _17891_ (
    .A(_6236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_6809_)
);

OR2X2 _17471_ (
    .A(_6388_),
    .B(_6395_),
    .Y(_6396_)
);

FILL FILL_0__17186_ (
);

AND2X2 _17051_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_5981_)
);

FILL FILL481080x350740 (
);

FILL FILL90440x54340 (
);

FILL FILL398240x360620 (
);

OR2X2 _9393_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_487_)
);

FILL FILL_0__10214_ (
);

AND2X2 _18676_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_7582_)
);

AND2X2 _18256_ (
    .A(_6289__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_7168_)
);

FILL FILL232560x291460 (
);

AND2X2 _13391_ (
    .A(_2925_),
    .B(_2927_),
    .Y(_2928_)
);

FILL FILL_0__19332_ (
);

FILL FILL253080x0 (
);

FILL FILL_0__11839_ (
);

OR2X2 _11704_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .B(_1718__bF$buf0),
    .Y(_1668_)
);

FILL FILL52440x311220 (
);

DFFSR _14596_ (
    .CLK(clk_bF$buf2),
    .D(_3738_[2]),
    .Q(\aluControl_1.inst [2]),
    .R(rst_bF$buf33),
    .S(vdd)
);

OR2X2 _14176_ (
    .A(MemToReg_bF$buf1),
    .B(ALUOut[11]),
    .Y(_3562_)
);

FILL FILL_0__15672_ (
);

FILL FILL471200x14820 (
);

AND2X2 _12909_ (
    .A(_2465_),
    .B(_2473_),
    .Y(_2474_)
);

FILL FILL286520x227240 (
);

FILL FILL_1_BUFX2_insert394 (
);

FILL FILL_1_BUFX2_insert396 (
);

FILL FILL_1_BUFX2_insert398 (
);

FILL FILL_1__17884_ (
);

FILL FILL_1__17464_ (
);

OR2X2 _10096_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .B(_860__bF$buf3),
    .Y(_856_)
);

FILL FILL240160x4940 (
);

OR2X2 _16742_ (
    .A(_5676_),
    .B(_5675_),
    .Y(_5677_)
);

FILL FILL_0__16457_ (
);

FILL FILL120840x158080 (
);

FILL FILL_0__16037_ (
);

AND2X2 _16322_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_5263_)
);

FILL FILL_0__11172_ (
);

OR2X2 _8664_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_121_)
);

FILL FILL203680x44460 (
);

AND2X2 _17947_ (
    .A(_6247__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_6864_)
);

OR2X2 _17527_ (
    .A(_6450_),
    .B(_6449_),
    .Y(_6451_)
);

OR2X2 _17107_ (
    .A(_6034_),
    .B(_6035_),
    .Y(_6036_)
);

FILL FILL_0__12797_ (
);

INVX1 _12662_ (
    .A(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2227_)
);

FILL FILL_0__12377_ (
);

AND2X2 _12242_ (
    .A(_1946_),
    .B(_1945_),
    .Y(_1917_[14])
);

FILL FILL_0__18603_ (
);

DFFSR _9869_ (
    .CLK(clk_bF$buf55),
    .D(_663_[26]),
    .Q(\datapath_1.regfile_1.regOut[11] [26]),
    .R(rst_bF$buf24),
    .S(vdd)
);

AND2X2 _9449_ (
    .A(_524_),
    .B(_523_),
    .Y(_465_[29])
);

AND2X2 _9029_ (
    .A(_304_),
    .B(_303_),
    .Y(_267_[18])
);

FILL FILL124640x266760 (
);

OR2X2 _13867_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [17]),
    .Y(_3311_)
);

AND2X2 _13447_ (
    .A(_2979_),
    .B(_2587_),
    .Y(_2980_)
);

AND2X2 _13027_ (
    .A(_2585_),
    .B(_2580_),
    .Y(_2586_)
);

FILL FILL_1__15530_ (
);

FILL FILL90440x345800 (
);

FILL FILL230280x340860 (
);

FILL FILL_0__14943_ (
);

FILL FILL_0__14523_ (
);

FILL FILL_0__14103_ (
);

FILL FILL261440x326040 (
);

FILL FILL452200x88920 (
);

AND2X2 _17280_ (
    .A(_6205_),
    .B(_6201_),
    .Y(_6206_)
);

FILL FILL_0__9909_ (
);

FILL FILL_0__15728_ (
);

FILL FILL_0__15308_ (
);

FILL FILL18240x29640 (
);

FILL FILL_0__10443_ (
);

FILL FILL_0__10023_ (
);

AND2X2 _18485_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_7394_)
);

NOR2X1 _18065_ (
    .A(_6310__bF$buf0),
    .B(_6979_),
    .Y(_6980_)
);

FILL FILL_1__12235_ (
);

FILL FILL_0__9662_ (
);

FILL FILL_0__11648_ (
);

DFFSR _11933_ (
    .CLK(clk_bF$buf89),
    .D(_1719_[26]),
    .Q(\datapath_1.regfile_1.regOut[27] [26]),
    .R(rst_bF$buf83),
    .S(vdd)
);

FILL FILL_0__11228_ (
);

AND2X2 _11513_ (
    .A(_1580_),
    .B(_1579_),
    .Y(_1521_[29])
);

FILL FILL300200x350740 (
);

FILL FILL46360x187720 (
);

FILL FILL_0__15481_ (
);

FILL FILL382280x256880 (
);

FILL FILL_0__15061_ (
);

FILL FILL82840x360620 (
);

FILL FILL299440x266760 (
);

FILL FILL63840x197600 (
);

XNOR2X1 _12718_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2283_)
);

FILL FILL_1_BUFX2_insert64 (
);

FILL FILL_1_BUFX2_insert66 (
);

FILL FILL_1_BUFX2_insert68 (
);

FILL FILL_0__16686_ (
);

AND2X2 _16971_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_5902_)
);

OR2X2 _16551_ (
    .A(_5485_),
    .B(_5488_),
    .Y(_5489_)
);

FILL FILL311600x44460 (
);

AND2X2 _16131_ (
    .A(_4160__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_5075_)
);

FILL FILL104120x44460 (
);

OR2X2 _8893_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .B(_266__bF$buf1),
    .Y(_234_)
);

OR2X2 _8473_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .B(_68__bF$buf3),
    .Y(_14_)
);

FILL FILL_1__13193_ (
);

OR2X2 _17756_ (
    .A(_6672_),
    .B(_6675_),
    .Y(_6676_)
);

AND2X2 _17336_ (
    .A(_6258_),
    .B(_6204_),
    .Y(_6262_)
);

OR2X2 _12891_ (
    .A(_2455_),
    .B(_2449_),
    .Y(_2456_)
);

AND2X2 _12471_ (
    .A(_2051_),
    .B(_2063_),
    .Y(_2064_)
);

DFFSR _12051_ (
    .CLK(clk_bF$buf51),
    .D(_1785_[15]),
    .Q(\datapath_1.regfile_1.regOut[28] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL413440x39520 (
);

FILL FILL449920x311220 (
);

FILL FILL_0__18832_ (
);

FILL FILL114000x158080 (
);

OR2X2 _9678_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_637_)
);

OR2X2 _9258_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_417_)
);

FILL FILL_0__8933_ (
);

FILL FILL_0__8513_ (
);

FILL FILL_0__10919_ (
);

FILL FILL_1_BUFX2_insert1154 (
);

AND2X2 _13676_ (
    .A(_3084__bF$buf4),
    .B(\datapath_1.PCJump [12]),
    .Y(_3159_)
);

OR2X2 _13256_ (
    .A(_2426_),
    .B(_2415_),
    .Y(_2801_)
);

FILL FILL_1_BUFX2_insert1156 (
);

FILL FILL_1_BUFX2_insert1158 (
);

FILL FILL473480x59280 (
);

FILL FILL370120x172900 (
);

FILL FILL_0__14332_ (
);

FILL FILL335160x335920 (
);

FILL FILL_0__15957_ (
);

FILL FILL_0__15537_ (
);

AND2X2 _15822_ (
    .A(_4167__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_4771_)
);

AND2X2 _15402_ (
    .A(_4197__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_4358_)
);

FILL FILL243200x4940 (
);

FILL FILL101080x148200 (
);

AND2X2 _18294_ (
    .A(_6302__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_7206_)
);

FILL FILL_0__19370_ (
);

FILL FILL433200x212420 (
);

FILL FILL_1__17749_ (
);

FILL FILL_1__17329_ (
);

OR2X2 _16607_ (
    .A(_5542_),
    .B(_5543_),
    .Y(_5544_)
);

FILL FILL_0__9891_ (
);

FILL FILL32680x143260 (
);

FILL FILL_0__11457_ (
);

OR2X2 _11742_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_1693_)
);

OR2X2 _11322_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_1473_)
);

OR2X2 _19499_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_8368_)
);

OR2X2 _19079_ (
    .A(_7977_),
    .B(_7978_),
    .Y(_7979_)
);

FILL FILL424080x316160 (
);

DFFSR _8949_ (
    .CLK(clk_bF$buf89),
    .D(_201_[9]),
    .Q(\datapath_1.regfile_1.regOut[4] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

OR2X2 _8529_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_51_)
);

FILL FILL_0__15290_ (
);

FILL FILL373920x44460 (
);

FILL FILL185440x316160 (
);

AND2X2 _12947_ (
    .A(_2510_),
    .B(_2497_),
    .Y(_2511_)
);

NOR2X1 _12527_ (
    .A(\control_1.reg_state.dout [2]),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2117_)
);

AND2X2 _12107_ (
    .A(_1876_),
    .B(_1875_),
    .Y(_1851_[12])
);

FILL FILL_1_BUFX2_insert774 (
);

FILL FILL_1_BUFX2_insert776 (
);

FILL FILL_1_BUFX2_insert778 (
);

FILL FILL281200x0 (
);

FILL FILL_0__13603_ (
);

FILL FILL440800x83980 (
);

OR2X2 _16780_ (
    .A(_5712_),
    .B(_5713_),
    .Y(_5714_)
);

FILL FILL186200x59280 (
);

FILL FILL_0__16075_ (
);

OR2X2 _16360_ (
    .A(_5300_),
    .B(_5293_),
    .Y(_5301_)
);

FILL FILL233320x83980 (
);

FILL FILL67640x237120 (
);

BUFX2 BUFX2_insert440 (
    .A(_1124_),
    .Y(_1124__bF$buf0)
);

BUFX2 BUFX2_insert441 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf4 )
);

BUFX2 BUFX2_insert442 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf3 )
);

BUFX2 BUFX2_insert443 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf2 )
);

BUFX2 BUFX2_insert444 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf1 )
);

AND2X2 _17985_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_6902_)
);

AND2X2 _17565_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_6488_)
);

BUFX2 BUFX2_insert445 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf0 )
);

FILL FILL453720x0 (
);

BUFX2 BUFX2_insert446 (
    .A(_1256_),
    .Y(_1256__bF$buf4)
);

OR2X2 _17145_ (
    .A(_6042_),
    .B(_6073_),
    .Y(_6074_)
);

BUFX2 BUFX2_insert447 (
    .A(_1256_),
    .Y(_1256__bF$buf3)
);

BUFX2 BUFX2_insert448 (
    .A(_1256_),
    .Y(_1256__bF$buf2)
);

BUFX2 BUFX2_insert449 (
    .A(_1256_),
    .Y(_1256__bF$buf1)
);

OR2X2 _12280_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_1982__bF$buf1),
    .Y(_1972_)
);

FILL FILL471960x148200 (
);

FILL FILL_0__18221_ (
);

FILL FILL370880x167960 (
);

DFFSR _9487_ (
    .CLK(clk_bF$buf57),
    .D(_465_[31]),
    .Q(\datapath_1.regfile_1.regOut[8] [31]),
    .R(rst_bF$buf81),
    .S(vdd)
);

OR2X2 _9067_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .B(_332__bF$buf4),
    .Y(_330_)
);

FILL FILL_1__11735_ (
);

FILL FILL_0__10728_ (
);

FILL FILL393680x251940 (
);

OR2X2 _13485_ (
    .A(RegDst),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_3013_)
);

AND2X2 _13065_ (
    .A(_2621_),
    .B(_2612_),
    .Y(_2622_)
);

FILL FILL_0__14561_ (
);

FILL FILL127680x182780 (
);

FILL FILL293360x345800 (
);

FILL FILL3800x143260 (
);

FILL FILL_0__9527_ (
);

FILL FILL_0__9107_ (
);

FILL FILL_1__16353_ (
);

OR2X2 _15631_ (
    .A(_4582_),
    .B(_4581_),
    .Y(_4583_)
);

NOR2X1 _15211_ (
    .A(_4144_),
    .B(_4140_),
    .Y(_4169_)
);

FILL FILL423320x167960 (
);

FILL FILL_0__10481_ (
);

FILL FILL335920x74100 (
);

FILL FILL150480x360620 (
);

FILL FILL_1__17978_ (
);

FILL FILL_1__12693_ (
);

OR2X2 _16836_ (
    .A(_5767_),
    .B(_5768_),
    .Y(_5769_)
);

OR2X2 _16416_ (
    .A(_5352_),
    .B(_5355_),
    .Y(_5356_)
);

FILL FILL_0__11686_ (
);

FILL FILL_0__9280_ (
);

OR2X2 _11971_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .B(_1850__bF$buf0),
    .Y(_1806_)
);

DFFSR _11551_ (
    .CLK(clk_bF$buf9),
    .D(_1521_[31]),
    .Q(\datapath_1.regfile_1.regOut[24] [31]),
    .R(rst_bF$buf23),
    .S(vdd)
);

OR2X2 _11131_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .B(_1388__bF$buf2),
    .Y(_1386_)
);

FILL FILL_0__17912_ (
);

OR2X2 _8758_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .B(_200__bF$buf4),
    .Y(_164_)
);

FILL FILL181640x14820 (
);

FILL FILL_1__13058_ (
);

FILL FILL285760x360620 (
);

OR2X2 _12756_ (
    .A(_2318_),
    .B(_2320_),
    .Y(_2321_)
);

OR2X2 _12336_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_1989_)
);

FILL FILL399760x108680 (
);

FILL FILL_0__13832_ (
);

FILL FILL404320x113620 (
);

FILL FILL415720x182780 (
);

FILL FILL11400x365560 (
);

AND2X2 _14902_ (
    .A(_3947_),
    .B(_3946_),
    .Y(_3936_[5])
);

OR2X2 _17794_ (
    .A(_6713_),
    .B(_6712_),
    .Y(_6714_)
);

AND2X2 _17374_ (
    .A(_6254_),
    .B(\datapath_1.PCJump_27_bF$buf0 ),
    .Y(_6300_)
);

FILL FILL_0__18870_ (
);

FILL FILL_0__18450_ (
);

FILL FILL15200x286520 (
);

FILL FILL_1__16829_ (
);

AND2X2 _9296_ (
    .A(_442_),
    .B(_441_),
    .Y(_399_[21])
);

FILL FILL_1__11124_ (
);

FILL FILL47120x74100 (
);

FILL FILL_0__8551_ (
);

FILL FILL_0__10957_ (
);

OR2X2 _10822_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .B(_1256__bF$buf1),
    .Y(_1220_)
);

FILL FILL_0__10537_ (
);

OR2X2 _10402_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .B(_1058__bF$buf0),
    .Y(_1000_)
);

OR2X2 _18999_ (
    .A(_7899_),
    .B(_7886_),
    .Y(_7900_)
);

FILL FILL383800x103740 (
);

OR2X2 _18579_ (
    .A(_7453_),
    .B(_7486_),
    .Y(_7487_)
);

FILL FILL66120x103740 (
);

AND2X2 _18159_ (
    .A(_6255__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_7073_)
);

FILL FILL29640x247000 (
);

XOR2X1 _13294_ (
    .A(_2219_),
    .B(_2210_),
    .Y(_2836_)
);

OR2X2 _19520_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_8382_)
);

FILL FILL_0__19235_ (
);

AND2X2 _19100_ (
    .A(_7999_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd1 [26])
);

FILL FILL_0__14370_ (
);

OR2X2 _11607_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_1623_)
);

FILL FILL283480x222300 (
);

OR2X2 _14499_ (
    .A(memoryOutData[0]),
    .B(_3803__bF$buf2),
    .Y(_3739_)
);

AND2X2 _14079_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3487_)
);

FILL FILL_1__16582_ (
);

AND2X2 _15860_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_4809_)
);

FILL FILL_0__15575_ (
);

FILL FILL_0__15155_ (
);

OR2X2 _15440_ (
    .A(_4391_),
    .B(_4394_),
    .Y(_4395_)
);

NOR2X1 _15020_ (
    .A(_4002_),
    .B(\datapath_1.a3 [1]),
    .Y(_4009_)
);

FILL FILL_0__10290_ (
);

FILL FILL3040x187720 (
);

FILL FILL505400x321100 (
);

AND2X2 _16645_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_5581_)
);

AND2X2 _16225_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_5168_)
);

FILL FILL_0__11495_ (
);

DFFSR _11780_ (
    .CLK(clk_bF$buf111),
    .D(_1653_[2]),
    .Q(\datapath_1.regfile_1.regOut[26] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

AND2X2 _11360_ (
    .A(_1498_),
    .B(_1497_),
    .Y(_1455_[21])
);

FILL FILL_0__11075_ (
);

FILL FILL_0__17721_ (
);

FILL FILL_0__17301_ (
);

AND2X2 _8987_ (
    .A(_276_),
    .B(_275_),
    .Y(_267_[4])
);

DFFSR _8567_ (
    .CLK(clk_bF$buf37),
    .D(_3_[14]),
    .Q(\datapath_1.regfile_1.regOut[1] [14]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_1__10815_ (
);

OR2X2 _12985_ (
    .A(_2157__bF$buf0),
    .B(_2545_),
    .Y(_2546_)
);

FILL FILL_1__19513_ (
);

AND2X2 _12565_ (
    .A(_2113_),
    .B(\control_1.op [1]),
    .Y(_2086_)
);

OR2X2 _12145_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .B(_1916__bF$buf4),
    .Y(_1902_)
);

FILL FILL_0__13641_ (
);

FILL FILL_0__13221_ (
);

FILL FILL448400x138320 (
);

FILL FILL_0__8607_ (
);

BUFX2 BUFX2_insert1000 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf4 )
);

BUFX2 BUFX2_insert1001 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf3 )
);

BUFX2 BUFX2_insert1002 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf2 )
);

BUFX2 BUFX2_insert1003 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf1 )
);

BUFX2 BUFX2_insert1004 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf0 )
);

BUFX2 BUFX2_insert1005 (
    .A(_3803_),
    .Y(_3803__bF$buf4)
);

BUFX2 BUFX2_insert1006 (
    .A(_3803_),
    .Y(_3803__bF$buf3)
);

BUFX2 BUFX2_insert1007 (
    .A(_3803_),
    .Y(_3803__bF$buf2)
);

BUFX2 BUFX2_insert1008 (
    .A(_3803_),
    .Y(_3803__bF$buf1)
);

BUFX2 BUFX2_insert1009 (
    .A(_3803_),
    .Y(_3803__bF$buf0)
);

FILL FILL_0__14846_ (
);

OR2X2 _14711_ (
    .A(vdd),
    .B(\datapath_1.a [28]),
    .Y(_3860_)
);

BUFX2 BUFX2_insert820 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf2 )
);

FILL FILL275880x103740 (
);

BUFX2 BUFX2_insert821 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf1 )
);

BUFX2 BUFX2_insert822 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf0 )
);

BUFX2 BUFX2_insert823 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf4 )
);

BUFX2 BUFX2_insert824 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf3 )
);

BUFX2 BUFX2_insert825 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf2 )
);

FILL FILL132240x133380 (
);

FILL FILL271320x74100 (
);

OR2X2 _17183_ (
    .A(_6110_),
    .B(_6109_),
    .Y(_6111_)
);

BUFX2 BUFX2_insert826 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf1 )
);

BUFX2 BUFX2_insert827 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf0 )
);

BUFX2 BUFX2_insert828 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf4 )
);

BUFX2 BUFX2_insert829 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf3 )
);

FILL FILL_1__16218_ (
);

FILL FILL70680x247000 (
);

AND2X2 _15916_ (
    .A(_4210__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_4864_)
);

FILL FILL205200x247000 (
);

FILL FILL_0__8780_ (
);

DFFSR _10631_ (
    .CLK(clk_bF$buf22),
    .D(_1059_[14]),
    .Q(\datapath_1.regfile_1.regOut[17] [14]),
    .R(rst_bF$buf7),
    .S(vdd)
);

FILL FILL_0__10346_ (
);

AND2X2 _10211_ (
    .A(_912_),
    .B(_911_),
    .Y(_861_[25])
);

OR2X2 _18388_ (
    .A(_7296_),
    .B(_7297_),
    .Y(_7298_)
);

FILL FILL_0__19464_ (
);

FILL FILL_0__19044_ (
);

FILL FILL_1__12138_ (
);

FILL FILL_0__9565_ (
);

OR2X2 _11836_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_1784__bF$buf3),
    .Y(_1736_)
);

DFFSR _11416_ (
    .CLK(clk_bF$buf81),
    .D(_1455_[25]),
    .Q(\datapath_1.regfile_1.regOut[23] [25]),
    .R(rst_bF$buf13),
    .S(vdd)
);

FILL FILL20520x29640 (
);

FILL FILL421040x19760 (
);

FILL FILL22800x360620 (
);

FILL FILL32680x306280 (
);

FILL FILL292600x98800 (
);

FILL FILL_0__16589_ (
);

AND2X2 _16874_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_5807_)
);

FILL FILL_0__16169_ (
);

AND2X2 _16454_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_5393_)
);

AND2X2 _16034_ (
    .A(_4154__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_4980_)
);

FILL FILL362520x350740 (
);

FILL FILL_0__17950_ (
);

FILL FILL_0__17110_ (
);

OR2X2 _8796_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_189_)
);

FILL FILL_1__10204_ (
);

AND2X2 _17659_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_6581_)
);

OR2X2 _17239_ (
    .A(_6162_),
    .B(_6165_),
    .Y(_6166_)
);

NAND2X1 _12794_ (
    .A(_2358_),
    .B(_2357_),
    .Y(_2359_)
);

AND2X2 _12374_ (
    .A(_2014_),
    .B(_2013_),
    .Y(_1983_[15])
);

FILL FILL_0__12089_ (
);

FILL FILL_0__18735_ (
);

FILL FILL_0__18315_ (
);

OR2X2 _18600_ (
    .A(_7505_),
    .B(_7506_),
    .Y(_7507_)
);

FILL FILL165680x286520 (
);

FILL FILL_0__13450_ (
);

FILL FILL_0__13030_ (
);

FILL FILL_1__11829_ (
);

FILL FILL296400x98800 (
);

FILL FILL_0__8416_ (
);

FILL FILL233320x207480 (
);

AND2X2 _13999_ (
    .A(_3352__bF$buf1),
    .B(\datapath_1.PCJump [11]),
    .Y(_3419_)
);

OR2X2 _13579_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.PCJump [30]),
    .Y(_3074_)
);

FILL FILL320720x212420 (
);

AOI21X1 _13159_ (
    .A(_2283_),
    .B(_2707_),
    .C(_2709_),
    .Y(_2710_)
);

FILL FILL502360x163020 (
);

FILL FILL357960x335920 (
);

FILL FILL_0__14655_ (
);

OR2X2 _14940_ (
    .A(\datapath_1.mux_pcsrc.dout [18]),
    .B(_4001__bF$buf1),
    .Y(_3973_)
);

OR2X2 _14520_ (
    .A(memoryOutData[7]),
    .B(_3803__bF$buf1),
    .Y(_3753_)
);

AND2X2 _14100_ (
    .A(_3344__bF$buf2),
    .B(gnd),
    .Y(_3505_)
);

FILL FILL323760x9880 (
);

FILL FILL176320x158080 (
);

FILL FILL_1__16867_ (
);

FILL FILL_1__16447_ (
);

FILL FILL303240x9880 (
);

AND2X2 _15725_ (
    .A(_4223__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_4676_)
);

OR2X2 _15305_ (
    .A(_4254_),
    .B(_4261_),
    .Y(_4262_)
);

FILL FILL_0__10575_ (
);

OR2X2 _10860_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_1245_)
);

FILL FILL_0__10155_ (
);

OR2X2 _10440_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_1025_)
);

OR2X2 _10020_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_805_)
);

OR2X2 _18197_ (
    .A(_7106_),
    .B(_7109_),
    .Y(_7110_)
);

FILL FILL82840x29640 (
);

FILL FILL235600x296400 (
);

FILL FILL_0__19273_ (
);

FILL FILL119320x64220 (
);

FILL FILL_0__9794_ (
);

FILL FILL_0__9374_ (
);

AND2X2 _11645_ (
    .A(_1648_),
    .B(_1647_),
    .Y(_1587_[30])
);

AND2X2 _11225_ (
    .A(_1428_),
    .B(_1427_),
    .Y(_1389_[19])
);

FILL FILL_0__12721_ (
);

FILL FILL297920x182780 (
);

FILL FILL_0__15193_ (
);

FILL FILL196080x34580 (
);

FILL FILL_1__14933_ (
);

FILL FILL_0__13926_ (
);

FILL FILL_0__13506_ (
);

FILL FILL488680x79040 (
);

OR2X2 _16683_ (
    .A(_5618_),
    .B(_5617_),
    .Y(_5619_)
);

FILL FILL_0__16398_ (
);

OR2X2 _16263_ (
    .A(_5204_),
    .B(_5203_),
    .Y(_5205_)
);

FILL FILL12920x103740 (
);

FILL FILL115520x261820 (
);

FILL FILL_1__10013_ (
);

AND2X2 _17888_ (
    .A(_6232__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_6806_)
);

AND2X2 _17468_ (
    .A(_6238__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_6393_)
);

OR2X2 _17048_ (
    .A(_5977_),
    .B(_5970_),
    .Y(_5978_)
);

DFFSR _12183_ (
    .CLK(clk_bF$buf110),
    .D(_1851_[18]),
    .Q(\datapath_1.regfile_1.regOut[29] [18]),
    .R(rst_bF$buf74),
    .S(vdd)
);

FILL FILL_1__19131_ (
);

FILL FILL12160x330980 (
);

FILL FILL_0__18964_ (
);

FILL FILL_0__18544_ (
);

FILL FILL_0__8645_ (
);

AND2X2 _10916_ (
    .A(_1262_),
    .B(_1261_),
    .Y(_1257_[2])
);

FILL FILL123880x375440 (
);

AND2X2 _13388_ (
    .A(_2923_),
    .B(_2924_),
    .Y(_2925_)
);

FILL FILL_1__15471_ (
);

FILL FILL_1__15051_ (
);

FILL FILL_0__19329_ (
);

FILL FILL_0__14884_ (
);

FILL FILL_0__14464_ (
);

FILL FILL_0__14044_ (
);

FILL FILL387600x321100 (
);

FILL FILL337440x172900 (
);

AND2X2 _15954_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_4901_)
);

FILL FILL_0__15669_ (
);

OR2X2 _15534_ (
    .A(_4486_),
    .B(_4487_),
    .Y(_4488_)
);

FILL FILL_0__15249_ (
);

AND2X2 _15114_ (
    .A(_4029_),
    .B(_4093_),
    .Y(\datapath_1.regfile_1.regEn [10])
);

FILL FILL_0__16610_ (
);

FILL FILL_0__19082_ (
);

OR2X2 _16739_ (
    .A(_5672_),
    .B(_5673_),
    .Y(_5674_)
);

AND2X2 _16319_ (
    .A(_4223__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_5260_)
);

OR2X2 _11874_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_1761_)
);

FILL FILL_0__11589_ (
);

OR2X2 _11454_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_1541_)
);

DFFSR _11034_ (
    .CLK(clk_bF$buf32),
    .D(_1257_[30]),
    .Q(\datapath_1.regfile_1.regOut[20] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL_0__17815_ (
);

FILL FILL_0__12950_ (
);

FILL FILL_0__12110_ (
);

FILL FILL253080x133380 (
);

DFFSR _9602_ (
    .CLK(clk_bF$buf8),
    .D(_531_[17]),
    .Q(\datapath_1.regfile_1.regOut[9] [17]),
    .R(rst_bF$buf73),
    .S(vdd)
);

OR2X2 _12659_ (
    .A(_2220_),
    .B(_2223_),
    .Y(_2224_)
);

AND2X2 _12239_ (
    .A(_1944_),
    .B(_1943_),
    .Y(_1917_[13])
);

FILL FILL_1__14322_ (
);

FILL FILL339720x108680 (
);

FILL FILL326040x247000 (
);

FILL FILL_0__13315_ (
);

OR2X2 _13600_ (
    .A(_3092_),
    .B(_3093_),
    .Y(_3094_)
);

FILL FILL411920x375440 (
);

FILL FILL_0_BUFX2_insert1160 (
);

FILL FILL_0_BUFX2_insert1161 (
);

FILL FILL_0_BUFX2_insert1162 (
);

FILL FILL_0_BUFX2_insert1163 (
);

AND2X2 _16492_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_5431_)
);

OR2X2 _16072_ (
    .A(_5016_),
    .B(_5013_),
    .Y(_5017_)
);

FILL FILL_0_BUFX2_insert1164 (
);

FILL FILL_0_BUFX2_insert1166 (
);

FILL FILL_0_BUFX2_insert1168 (
);

FILL FILL_1__15947_ (
);

OR2X2 _14805_ (
    .A(\datapath_1.rd2 [16]),
    .B(_3935__bF$buf0),
    .Y(_3903_)
);

FILL FILL159600x286520 (
);

OR2X2 _17697_ (
    .A(_6617_),
    .B(_6616_),
    .Y(_6618_)
);

AND2X2 _17277_ (
    .A(_6202_),
    .B(\datapath_1.PCJump [23]),
    .Y(_6203_)
);

FILL FILL88160x143260 (
);

FILL FILL_0__18353_ (
);

DFFSR _9199_ (
    .CLK(clk_bF$buf69),
    .D(_333_[1]),
    .Q(\datapath_1.regfile_1.regOut[6] [1]),
    .R(rst_bF$buf76),
    .S(vdd)
);

FILL FILL_1__11867_ (
);

FILL FILL_0__8454_ (
);

OR2X2 _10725_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_1175_)
);

OR2X2 _10305_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_955_)
);

AND2X2 _13197_ (
    .A(_2745_),
    .B(_2443_),
    .Y(_2746_)
);

FILL FILL377720x276640 (
);

OR2X2 _19423_ (
    .A(_8286_),
    .B(_8317_),
    .Y(_8318_)
);

FILL FILL_0__19138_ (
);

OR2X2 _19003_ (
    .A(_7902_),
    .B(_7903_),
    .Y(_7904_)
);

FILL FILL_0__14693_ (
);

FILL FILL_0__14273_ (
);

FILL FILL464360x187720 (
);

FILL FILL_0__9659_ (
);

FILL FILL_0__9239_ (
);

FILL FILL_0__15898_ (
);

FILL FILL234840x291460 (
);

OR2X2 _15763_ (
    .A(_4711_),
    .B(_4712_),
    .Y(_4713_)
);

FILL FILL_0__15058_ (
);

OR2X2 _15343_ (
    .A(_4296_),
    .B(_4299_),
    .Y(_4300_)
);

FILL FILL153520x227240 (
);

FILL FILL302480x29640 (
);

FILL FILL_1__8615_ (
);

FILL FILL31920x227240 (
);

OR2X2 _16968_ (
    .A(_5898_),
    .B(_5895_),
    .Y(_5899_)
);

AND2X2 _16548_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_5486_)
);

OR2X2 _16128_ (
    .A(_5071_),
    .B(_5070_),
    .Y(_5072_)
);

FILL FILL_1__18631_ (
);

OR2X2 _11683_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(_1718__bF$buf4),
    .Y(_1654_)
);

FILL FILL_1__18211_ (
);

DFFSR _11263_ (
    .CLK(clk_bF$buf43),
    .D(_1389_[1]),
    .Q(\datapath_1.regfile_1.regOut[22] [1]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL_0__17204_ (
);

FILL FILL361000x177840 (
);

OR2X2 _9831_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_719_)
);

OR2X2 _9411_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_499_)
);

NOR2X1 _12888_ (
    .A(_2282_),
    .B(_2283_),
    .Y(_2453_)
);

AND2X2 _12468_ (
    .A(_2060_),
    .B(\aluControl_1.inst [1]),
    .Y(_2061_)
);

DFFSR _12048_ (
    .CLK(clk_bF$buf93),
    .D(_1785_[12]),
    .Q(\datapath_1.regfile_1.regOut[28] [12]),
    .R(rst_bF$buf41),
    .S(vdd)
);

FILL FILL_0__18829_ (
);

FILL FILL_0__18409_ (
);

FILL FILL_0__13544_ (
);

FILL FILL433960x44460 (
);

FILL FILL471200x88920 (
);

FILL FILL_1__15336_ (
);

FILL FILL17480x14820 (
);

FILL FILL505400x281580 (
);

DFFSR _14614_ (
    .CLK(clk_bF$buf40),
    .D(_3738_[20]),
    .Q(\datapath_1.PCJump [22]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL_0__14329_ (
);

AND2X2 _17086_ (
    .A(_4187__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_6015_)
);

FILL FILL_0__18582_ (
);

FILL FILL_0__18162_ (
);

FILL FILL132240x247000 (
);

FILL FILL281200x153140 (
);

FILL FILL_1__11256_ (
);

AND2X2 _15819_ (
    .A(_4135__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_4768_)
);

FILL FILL126920x266760 (
);

OR2X2 _10954_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .B(_1322__bF$buf1),
    .Y(_1288_)
);

FILL FILL_0__10669_ (
);

OR2X2 _10534_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .B(_1124__bF$buf2),
    .Y(_1068_)
);

DFFSR _10114_ (
    .CLK(clk_bF$buf13),
    .D(_795_[13]),
    .Q(\datapath_1.regfile_1.regOut[13] [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

FILL FILL318440x355680 (
);

AND2X2 _19232_ (
    .A(_6293__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_8129_)
);

FILL FILL164160x222300 (
);

FILL FILL_0__14082_ (
);

OR2X2 _11739_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_1691_)
);

FILL FILL_0__9048_ (
);

OR2X2 _11319_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_1471_)
);

FILL FILL_1__13822_ (
);

FILL FILL_0__12815_ (
);

FILL FILL264480x0 (
);

OR2X2 _15992_ (
    .A(_4938_),
    .B(_4923_),
    .Y(_4939_)
);

FILL FILL_0__15287_ (
);

AND2X2 _15572_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_4525_)
);

AND2X2 _15152_ (
    .A(_4116_),
    .B(_4008_),
    .Y(_4117_)
);

FILL FILL253840x271700 (
);

FILL FILL_1__8424_ (
);

FILL FILL330600x44460 (
);

FILL FILL497040x98800 (
);

FILL FILL505400x54340 (
);

FILL FILL454480x251940 (
);

OR2X2 _16777_ (
    .A(_5703_),
    .B(_5710_),
    .Y(_5711_)
);

AND2X2 _16357_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_5298_)
);

FILL FILL_1__18860_ (
);

AND2X2 _11492_ (
    .A(_1566_),
    .B(_1565_),
    .Y(_1521_[22])
);

AND2X2 _11072_ (
    .A(_1346_),
    .B(_1345_),
    .Y(_1323_[11])
);

FILL FILL_1__9629_ (
);

FILL FILL48640x187720 (
);

FILL FILL_0__17853_ (
);

FILL FILL_0__17433_ (
);

DFFSR _8699_ (
    .CLK(clk_bF$buf8),
    .D(_69_[17]),
    .Q(\datapath_1.regfile_1.regOut[2] [17]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL_1__10947_ (
);

FILL FILL133000x251940 (
);

FILL FILL458280x172900 (
);

OR2X2 _9640_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_662__bF$buf1),
    .Y(_612_)
);

DFFSR _9220_ (
    .CLK(clk_bF$buf87),
    .D(_333_[22]),
    .Q(\datapath_1.regfile_1.regOut[6] [22]),
    .R(rst_bF$buf2),
    .S(vdd)
);

NAND2X1 _12697_ (
    .A(_2260_),
    .B(_2261_),
    .Y(_2262_)
);

OR2X2 _12277_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_1982__bF$buf0),
    .Y(_1970_)
);

FILL FILL230280x202540 (
);

FILL FILL_1__14780_ (
);

FILL FILL_0__18638_ (
);

AND2X2 _18923_ (
    .A(_6250__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_7825_)
);

FILL FILL_0__18218_ (
);

OR2X2 _18503_ (
    .A(_7411_),
    .B(_7408_),
    .Y(_7412_)
);

FILL FILL_0__13773_ (
);

FILL FILL_0__8739_ (
);

FILL FILL15200x172900 (
);

FILL FILL416480x24700 (
);

FILL FILL141360x365560 (
);

FILL FILL329840x123500 (
);

FILL FILL_1__15565_ (
);

FILL FILL35720x49400 (
);

FILL FILL25080x118560 (
);

FILL FILL_0__14978_ (
);

OR2X2 _14843_ (
    .A(vdd),
    .B(_2_[29]),
    .Y(_3928_)
);

FILL FILL_0__14138_ (
);

OR2X2 _14423_ (
    .A(vdd),
    .B(\datapath_1.Data [18]),
    .Y(_3708_)
);

AND2X2 _14003_ (
    .A(_3347__bF$buf0),
    .B(\datapath_1.PCJump [14]),
    .Y(_3422_)
);

FILL FILL433200x4940 (
);

FILL FILL145160x286520 (
);

FILL FILL_0__18391_ (
);

FILL FILL_1__11065_ (
);

OR2X2 _15628_ (
    .A(_4578_),
    .B(_4579_),
    .Y(_4580_)
);

AND2X2 _15208_ (
    .A(_4139_),
    .B(_4165_),
    .Y(_4166_)
);

FILL FILL_0__8492_ (
);

FILL FILL_0__10478_ (
);

FILL FILL_1__17711_ (
);

DFFSR _10763_ (
    .CLK(clk_bF$buf76),
    .D(_1125_[17]),
    .Q(\datapath_1.regfile_1.regOut[18] [17]),
    .R(rst_bF$buf112),
    .S(vdd)
);

AND2X2 _10343_ (
    .A(_980_),
    .B(_979_),
    .Y(_927_[26])
);

FILL FILL_0__10058_ (
);

FILL FILL477280x158080 (
);

FILL FILL196080x103740 (
);

FILL FILL327560x197600 (
);

FILL FILL_0__16704_ (
);

FILL FILL_0__19176_ (
);

OR2X2 _19461_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8343_)
);

OR2X2 _19041_ (
    .A(_7940_),
    .B(_7939_),
    .Y(_7941_)
);

OR2X2 _8911_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .B(_266__bF$buf4),
    .Y(_246_)
);

FILL FILL363280x276640 (
);

FILL FILL_0__9697_ (
);

OR2X2 _11968_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .B(_1850__bF$buf3),
    .Y(_1804_)
);

DFFSR _11548_ (
    .CLK(clk_bF$buf84),
    .D(_1521_[28]),
    .Q(\datapath_1.regfile_1.regOut[24] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

OR2X2 _11128_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_1388__bF$buf3),
    .Y(_1384_)
);

FILL FILL_0__17909_ (
);

FILL FILL_0__12624_ (
);

FILL FILL_0__12204_ (
);

FILL FILL103360x148200 (
);

FILL FILL63080x286520 (
);

FILL FILL386080x360620 (
);

FILL FILL_0__15096_ (
);

AND2X2 _15381_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_4337_)
);

FILL FILL_0__13409_ (
);

AND2X2 _16586_ (
    .A(_4203__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_5523_)
);

OR2X2 _16166_ (
    .A(_5109_),
    .B(_5108_),
    .Y(_5110_)
);

FILL FILL426360x316160 (
);

FILL FILL_1__9018_ (
);

FILL FILL_0__17662_ (
);

FILL FILL391400x158080 (
);

FILL FILL21280x148200 (
);

FILL FILL344280x222300 (
);

AND2X2 _12086_ (
    .A(_1862_),
    .B(_1861_),
    .Y(_1851_[5])
);

FILL FILL_0__18867_ (
);

AND2X2 _18732_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_7637_)
);

AND2X2 _18312_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_7224_)
);

FILL FILL_0__18027_ (
);

FILL FILL_0__13582_ (
);

FILL FILL_0__13162_ (
);

OR2X2 _10819_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_1256__bF$buf1),
    .Y(_1218_)
);

FILL FILL120080x74100 (
);

FILL FILL85120x0 (
);

OR2X2 _19517_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_8380_)
);

FILL FILL_0__14787_ (
);

OR2X2 _14652_ (
    .A(\datapath_1.rd1 [8]),
    .B(_3869__bF$buf2),
    .Y(_3821_)
);

AND2X2 _14232_ (
    .A(_3599_),
    .B(_3598_),
    .Y(\datapath_1.mux_wd3.dout [29])
);

FILL FILL501600x98800 (
);

FILL FILL278160x335920 (
);

AND2X2 _15857_ (
    .A(_4239__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_4806_)
);

AND2X2 _15437_ (
    .A(_4234__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_4392_)
);

NAND2X1 _15017_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_4006_)
);

OR2X2 _10992_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_1313_)
);

FILL FILL_0__10287_ (
);

OR2X2 _10572_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_1093_)
);

FILL FILL_1__17100_ (
);

OR2X2 _10152_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_873_)
);

FILL FILL496280x138320 (
);

FILL FILL_0__16933_ (
);

FILL FILL129960x182780 (
);

FILL FILL462080x93860 (
);

AND2X2 _19270_ (
    .A(_6315__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_8167_)
);

AND2X2 _8720_ (
    .A(_138_),
    .B(_137_),
    .Y(_135_[1])
);

FILL FILL_1__18725_ (
);

AND2X2 _11777_ (
    .A(_1716_),
    .B(_1715_),
    .Y(_1653_[31])
);

AND2X2 _11357_ (
    .A(_1496_),
    .B(_1495_),
    .Y(_1455_[20])
);

FILL FILL_1__13440_ (
);

FILL FILL_0__17718_ (
);

FILL FILL308560x370500 (
);

FILL FILL376200x212420 (
);

OR2X2 _15190_ (
    .A(_4143_),
    .B(_4147_),
    .Y(_4148_)
);

OR2X2 _9925_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .B(_794__bF$buf3),
    .Y(_762_)
);

OR2X2 _9505_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_596__bF$buf3),
    .Y(_542_)
);

FILL FILL484880x232180 (
);

FILL FILL17480x271700 (
);

OR2X2 _13923_ (
    .A(_3353_),
    .B(_3351_),
    .Y(_3354_)
);

FILL FILL_0__13638_ (
);

AND2X2 _13503_ (
    .A(_3023_),
    .B(_3022_),
    .Y(_1_[4])
);

FILL FILL87400x291460 (
);

AND2X2 _16395_ (
    .A(_4130__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_5335_)
);

FILL FILL_0__17471_ (
);

FILL FILL_0__17051_ (
);

FILL FILL488680x153140 (
);

FILL FILL_1__10565_ (
);

OR2X2 _14708_ (
    .A(vdd),
    .B(\datapath_1.a [27]),
    .Y(_3858_)
);

BUFX2 BUFX2_insert790 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf2 )
);

BUFX2 BUFX2_insert791 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf1 )
);

BUFX2 BUFX2_insert792 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf0 )
);

BUFX2 BUFX2_insert793 (
    .A(_4236_),
    .Y(_4236__bF$buf4)
);

BUFX2 BUFX2_insert794 (
    .A(_4236_),
    .Y(_4236__bF$buf3)
);

BUFX2 BUFX2_insert795 (
    .A(_4236_),
    .Y(_4236__bF$buf2)
);

BUFX2 BUFX2_insert796 (
    .A(_4236_),
    .Y(_4236__bF$buf1)
);

BUFX2 BUFX2_insert797 (
    .A(_4236_),
    .Y(_4236__bF$buf0)
);

BUFX2 BUFX2_insert798 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf4 )
);

BUFX2 BUFX2_insert799 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf3 )
);

FILL FILL28120x143260 (
);

FILL FILL319200x108680 (
);

FILL FILL406600x113620 (
);

FILL FILL_0__18676_ (
);

OR2X2 _18961_ (
    .A(_7861_),
    .B(_7862_),
    .Y(_7863_)
);

FILL FILL_0__18256_ (
);

AND2X2 _18541_ (
    .A(_6264__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_7449_)
);

OR2X2 _18121_ (
    .A(_7035_),
    .B(_7028_),
    .Y(_7036_)
);

FILL FILL302480x311220 (
);

FILL FILL_0__13391_ (
);

FILL FILL45600x153140 (
);

DFFSR _10628_ (
    .CLK(clk_bF$buf73),
    .D(_1059_[11]),
    .Q(\datapath_1.regfile_1.regOut[17] [11]),
    .R(rst_bF$buf39),
    .S(vdd)
);

AND2X2 _10208_ (
    .A(_910_),
    .B(_909_),
    .Y(_861_[24])
);

AND2X2 _19326_ (
    .A(_6282__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_8222_)
);

DFFSR _14881_ (
    .CLK(clk_bF$buf40),
    .D(_3870_[29]),
    .Q(_2_[29]),
    .R(rst_bF$buf63),
    .S(vdd)
);

AND2X2 _14461_ (
    .A(_3733_),
    .B(_3732_),
    .Y(_3672_[30])
);

AND2X2 _14041_ (
    .A(_3352__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3455_)
);

FILL FILL_1__13916_ (
);

FILL FILL_0__12909_ (
);

FILL FILL_1__16388_ (
);

FILL FILL245480x128440 (
);

OR2X2 _15666_ (
    .A(_4616_),
    .B(_4617_),
    .Y(_4618_)
);

AND2X2 _15246_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_4204_)
);

FILL FILL418760x148200 (
);

FILL FILL440040x266760 (
);

DFFSR _10381_ (
    .CLK(clk_bF$buf101),
    .D(_927_[22]),
    .Q(\datapath_1.regfile_1.regOut[15] [22]),
    .R(rst_bF$buf54),
    .S(vdd)
);

FILL FILL_0__10096_ (
);

FILL FILL_1__8518_ (
);

FILL FILL_0__16322_ (
);

FILL FILL243960x296400 (
);

FILL FILL285760x222300 (
);

OR2X2 _11586_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_1609_)
);

INVX2 _11166_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .Y(_1454_)
);

FILL FILL_0__17947_ (
);

FILL FILL_0__17527_ (
);

AND2X2 _17812_ (
    .A(_6216__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_6731_)
);

FILL FILL_0__12662_ (
);

FILL FILL389120x251940 (
);

DFFSR _9734_ (
    .CLK(clk_bF$buf95),
    .D(_597_[20]),
    .Q(\datapath_1.regfile_1.regOut[10] [20]),
    .R(rst_bF$buf30),
    .S(vdd)
);

AND2X2 _9314_ (
    .A(_454_),
    .B(_453_),
    .Y(_399_[27])
);

FILL FILL_1__14454_ (
);

FILL FILL_0__13867_ (
);

FILL FILL_0__13447_ (
);

AND2X2 _13732_ (
    .A(_3084__bF$buf2),
    .B(\datapath_1.PCJump [20]),
    .Y(_3207_)
);

FILL FILL_0__13027_ (
);

INVX1 _13312_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .Y(_2853_)
);

FILL FILL215840x54340 (
);

FILL FILL_0__17280_ (
);

OR2X2 _14937_ (
    .A(\datapath_1.mux_pcsrc.dout [17]),
    .B(_4001__bF$buf0),
    .Y(_3971_)
);

OR2X2 _14517_ (
    .A(memoryOutData[6]),
    .B(_3803__bF$buf0),
    .Y(_3751_)
);

FILL FILL_1__19072_ (
);

FILL FILL47120x123500 (
);

OR2X2 _18770_ (
    .A(_7671_),
    .B(_7674_),
    .Y(_7675_)
);

OR2X2 _18350_ (
    .A(_7247_),
    .B(_7260_),
    .Y(_7261_)
);

FILL FILL66880x44460 (
);

FILL FILL_1__11999_ (
);

OR2X2 _10857_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_1243_)
);

OR2X2 _10437_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_1023_)
);

OR2X2 _10017_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_803_)
);

FILL FILL_1__12940_ (
);

FILL FILL219640x54340 (
);

FILL FILL486400x217360 (
);

FILL FILL22800x79040 (
);

INVX1 _19555_ (
    .A(ALUZero),
    .Y(_8386_)
);

AND2X2 _19135_ (
    .A(_6315__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_8034_)
);

FILL FILL111720x83980 (
);

OR2X2 _14690_ (
    .A(vdd),
    .B(\datapath_1.a [21]),
    .Y(_3846_)
);

OR2X2 _14270_ (
    .A(vdd),
    .B(ALUOut[10]),
    .Y(_3626_)
);

FILL FILL499320x163020 (
);

FILL FILL467400x375440 (
);

FILL FILL_1__13305_ (
);

FILL FILL72960x247000 (
);

OR2X2 _15895_ (
    .A(_4839_),
    .B(_4842_),
    .Y(_4843_)
);

AND2X2 _15475_ (
    .A(_4228__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_4430_)
);

NAND2X1 _15055_ (
    .A(_4024_),
    .B(_4030_),
    .Y(_4044_)
);

AND2X2 _10190_ (
    .A(_898_),
    .B(_897_),
    .Y(_861_[18])
);

FILL FILL_0__16971_ (
);

FILL FILL_0__16551_ (
);

FILL FILL203680x217360 (
);

FILL FILL_0__16131_ (
);

FILL FILL467400x19760 (
);

FILL FILL430920x103740 (
);

DFFSR _11395_ (
    .CLK(clk_bF$buf73),
    .D(_1455_[4]),
    .Q(\datapath_1.regfile_1.regOut[23] [4]),
    .R(rst_bF$buf39),
    .S(vdd)
);

FILL FILL_0__17756_ (
);

OR2X2 _17621_ (
    .A(_6534_),
    .B(_6542_),
    .Y(_6543_)
);

FILL FILL_0__17336_ (
);

AND2X2 _17201_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_6129_)
);

FILL FILL_0__12891_ (
);

FILL FILL430160x330980 (
);

OR2X2 _9963_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_787_)
);

OR2X2 _9543_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_567_)
);

OR2X2 _9123_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [7]),
    .Y(_347_)
);

FILL FILL338960x217360 (
);

FILL FILL_1__14263_ (
);

AND2X2 _18826_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_7730_)
);

FILL FILL_0_BUFX2_insert431 (
);

AND2X2 _18406_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_7316_)
);

FILL FILL_0_BUFX2_insert433 (
);

AND2X2 _13961_ (
    .A(_3347__bF$buf1),
    .B(\datapath_1.PCJump [8]),
    .Y(_3386_)
);

FILL FILL_0__13256_ (
);

FILL FILL_0_BUFX2_insert435 (
);

OR2X2 _13541_ (
    .A(ALUOut[17]),
    .B(_3079__bF$buf1),
    .Y(_3049_)
);

AOI21X1 _13121_ (
    .A(_2280_),
    .B(_2504_),
    .C(_2673_),
    .Y(_2674_)
);

FILL FILL_0_BUFX2_insert437 (
);

FILL FILL319960x375440 (
);

FILL FILL_0_BUFX2_insert438 (
);

FILL FILL_0_BUFX2_insert439 (
);

FILL FILL256880x123500 (
);

FILL FILL137560x93860 (
);

FILL FILL321480x93860 (
);

FILL FILL459800x256880 (
);

FILL FILL_1__15888_ (
);

FILL FILL186960x128440 (
);

DFFSR _14746_ (
    .CLK(clk_bF$buf94),
    .D(_3804_[23]),
    .Q(\datapath_1.a [23]),
    .R(rst_bF$buf61),
    .S(vdd)
);

AND2X2 _14326_ (
    .A(_3663_),
    .B(_3662_),
    .Y(_3606_[28])
);

FILL FILL_0__15822_ (
);

FILL FILL_0__15402_ (
);

FILL FILL_0__18294_ (
);

OR2X2 _10666_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_1190__bF$buf4),
    .Y(_1136_)
);

DFFSR _10246_ (
    .CLK(clk_bF$buf8),
    .D(_861_[16]),
    .Q(\datapath_1.regfile_1.regOut[14] [16]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL417240x158080 (
);

FILL FILL504640x163020 (
);

FILL FILL248520x153140 (
);

FILL FILL499320x256880 (
);

FILL FILL_0__11742_ (
);

FILL FILL_0__19499_ (
);

AND2X2 _19364_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_8259_)
);

FILL FILL313880x316160 (
);

DFFSR _8814_ (
    .CLK(clk_bF$buf10),
    .D(_135_[3]),
    .Q(\datapath_1.regfile_1.regOut[3] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL284240x232180 (
);

FILL FILL_1__13954_ (
);

INVX1 _12812_ (
    .A(_2159_),
    .Y(_2377_)
);

FILL FILL_0__12527_ (
);

FILL FILL_0__12107_ (
);

FILL FILL389880x197600 (
);

AND2X2 _15284_ (
    .A(_4241__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_4242_)
);

FILL FILL_0__16780_ (
);

AND2X2 _16489_ (
    .A(_4158__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_5428_)
);

AND2X2 _16069_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_5014_)
);

FILL FILL438520x276640 (
);

FILL FILL96520x158080 (
);

FILL FILL174040x271700 (
);

FILL FILL_1__18152_ (
);

FILL FILL_0__17985_ (
);

AND2X2 _17850_ (
    .A(_6287__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_6769_)
);

OR2X2 _17430_ (
    .A(_6352_),
    .B(_6354_),
    .Y(_6355_)
);

FILL FILL_0__17145_ (
);

OR2X2 _17010_ (
    .A(_5939_),
    .B(_5940_),
    .Y(_5941_)
);

FILL FILL_0__12280_ (
);

FILL FILL_1__10659_ (
);

FILL FILL92720x83980 (
);

OR2X2 _9772_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .B(_728__bF$buf4),
    .Y(_680_)
);

DFFSR _9352_ (
    .CLK(clk_bF$buf81),
    .D(_399_[25]),
    .Q(\datapath_1.regfile_1.regOut[7] [25]),
    .R(rst_bF$buf101),
    .S(vdd)
);

AND2X2 _18635_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_7542_)
);

AND2X2 _18215_ (
    .A(_6264__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_7128_)
);

FILL FILL_0__13485_ (
);

AND2X2 _13770_ (
    .A(_3089__bF$buf2),
    .B(gnd),
    .Y(_3240_)
);

FILL FILL_0__13065_ (
);

INVX1 _13350_ (
    .A(_2889_),
    .Y(\datapath_1.ALUResult [6])
);

FILL FILL200640x251940 (
);

FILL FILL_1__12805_ (
);

FILL FILL_0__9812_ (
);

OR2X2 _14975_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.PCJump [30]),
    .Y(_3996_)
);

OR2X2 _14555_ (
    .A(IRWrite_bF$buf0),
    .B(\datapath_1.PCJump [21]),
    .Y(_3776_)
);

AND2X2 _14135_ (
    .A(_3344__bF$buf1),
    .B(gnd),
    .Y(_3535_)
);

FILL FILL419520x222300 (
);

FILL FILL186200x9880 (
);

FILL FILL504640x256880 (
);

DFFSR _10895_ (
    .CLK(clk_bF$buf9),
    .D(_1191_[20]),
    .Q(\datapath_1.regfile_1.regOut[19] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

FILL FILL_1__17843_ (
);

AND2X2 _10475_ (
    .A(_1048_),
    .B(_1047_),
    .Y(_993_[27])
);

AND2X2 _10055_ (
    .A(_828_),
    .B(_827_),
    .Y(_795_[16])
);

FILL FILL49400x237120 (
);

FILL FILL_0__16836_ (
);

OR2X2 _16701_ (
    .A(_5635_),
    .B(_5634_),
    .Y(_5636_)
);

FILL FILL_0__16416_ (
);

FILL FILL_0__11971_ (
);

FILL FILL_0__11131_ (
);

FILL FILL44080x192660 (
);

AND2X2 _19173_ (
    .A(_6229__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_8071_)
);

OR2X2 _8623_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .B(_134__bF$buf1),
    .Y(_94_)
);

OR2X2 _17906_ (
    .A(_6822_),
    .B(_6823_),
    .Y(_6824_)
);

FILL FILL_0__12756_ (
);

XNOR2X1 _12621_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2186_)
);

FILL FILL_0__12336_ (
);

OR2X2 _12201_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_1919_)
);

AND2X2 _15093_ (
    .A(_4070_),
    .B(_4076_),
    .Y(_4077_)
);

OR2X2 _9828_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_717_)
);

OR2X2 _9408_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_497_)
);

FILL FILL_1__14128_ (
);

OR2X2 _13826_ (
    .A(\datapath_1.a [3]),
    .B(_3342__bF$buf1),
    .Y(_3284_)
);

OR2X2 _13406_ (
    .A(_2930_),
    .B(_2501_),
    .Y(_2942_)
);

FILL FILL414200x192660 (
);

AND2X2 _16298_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_5240_)
);

FILL FILL_0__14902_ (
);

FILL FILL487920x167960 (
);

FILL FILL255360x133380 (
);

FILL FILL_0__17794_ (
);

FILL FILL_0__17374_ (
);

FILL FILL411160x237120 (
);

AND2X2 _9581_ (
    .A(_592_),
    .B(_591_),
    .Y(_531_[30])
);

AND2X2 _9161_ (
    .A(_372_),
    .B(_371_),
    .Y(_333_[19])
);

FILL FILL_1__19166_ (
);

FILL FILL_0__10822_ (
);

FILL FILL_0__18999_ (
);

AND2X2 _18864_ (
    .A(_6321__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_7767_)
);

FILL FILL_0__18159_ (
);

FILL FILL_0_BUFX2_insert811 (
);

OR2X2 _18444_ (
    .A(_7353_),
    .B(_7352_),
    .Y(_7354_)
);

FILL FILL314640x271700 (
);

OR2X2 _18024_ (
    .A(_6939_),
    .B(_6926_),
    .Y(_6940_)
);

FILL FILL_0_BUFX2_insert813 (
);

FILL FILL_0_BUFX2_insert815 (
);

FILL FILL57760x34580 (
);

FILL FILL_0_BUFX2_insert817 (
);

FILL FILL_0_BUFX2_insert818 (
);

FILL FILL_0_BUFX2_insert819 (
);

FILL FILL_0__19100_ (
);

FILL FILL350360x350740 (
);

FILL FILL_0__9621_ (
);

FILL FILL_0__11607_ (
);

OR2X2 _19229_ (
    .A(_8092_),
    .B(_8126_),
    .Y(_8127_)
);

OR2X2 _14784_ (
    .A(\datapath_1.rd2 [9]),
    .B(_3935__bF$buf1),
    .Y(_3889_)
);

FILL FILL_0__14079_ (
);

DFFSR _14364_ (
    .CLK(clk_bF$buf50),
    .D(_3606_[28]),
    .Q(ALUOut[28]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL_0__15440_ (
);

FILL FILL_0__15020_ (
);

FILL FILL449920x271700 (
);

OR2X2 _15989_ (
    .A(_4935_),
    .B(_4934_),
    .Y(_4936_)
);

AND2X2 _15569_ (
    .A(_4151__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_4522_)
);

AND2X2 _15149_ (
    .A(_4115_),
    .B(_4112_),
    .Y(\datapath_1.regfile_1.regEn [23])
);

OR2X2 _10284_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_941_)
);

FILL FILL_0__16645_ (
);

AND2X2 _16930_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_5862_)
);

AND2X2 _16510_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_5448_)
);

FILL FILL_0__16225_ (
);

FILL FILL485640x350740 (
);

FILL FILL_0__11360_ (
);

FILL FILL293360x167960 (
);

FILL FILL79800x286520 (
);

AND2X2 _8852_ (
    .A(_206_),
    .B(_205_),
    .Y(_201_[2])
);

BUFX2 _8432_ (
    .A(_2_[8]),
    .Y(memoryWriteData[8])
);

FILL FILL34200x19760 (
);

AND2X2 _11489_ (
    .A(_1564_),
    .B(_1563_),
    .Y(_1521_[21])
);

AND2X2 _11069_ (
    .A(_1344_),
    .B(_1343_),
    .Y(_1323_[10])
);

FILL FILL_1__18017_ (
);

FILL FILL119320x375440 (
);

OR2X2 _17715_ (
    .A(_6632_),
    .B(_6635_),
    .Y(_6636_)
);

FILL FILL_0__12985_ (
);

AND2X2 _12850_ (
    .A(_2405_),
    .B(_2414_),
    .Y(_2415_)
);

FILL FILL_0__12145_ (
);

DFFSR _12430_ (
    .CLK(clk_bF$buf66),
    .D(_1983_[7]),
    .Q(\datapath_1.regfile_1.regOut[31] [7]),
    .R(rst_bF$buf80),
    .S(vdd)
);

OR2X2 _12010_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .B(_1850__bF$buf4),
    .Y(_1832_)
);

FILL FILL185440x0 (
);

OR2X2 _9637_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .B(_662__bF$buf1),
    .Y(_610_)
);

DFFSR _9217_ (
    .CLK(clk_bF$buf69),
    .D(_333_[19]),
    .Q(\datapath_1.regfile_1.regOut[6] [19]),
    .R(rst_bF$buf13),
    .S(vdd)
);

OR2X2 _13635_ (
    .A(_3122_),
    .B(_3123_),
    .Y(_3124_)
);

AND2X2 _13215_ (
    .A(_2762_),
    .B(_2754_),
    .Y(_2763_)
);

FILL FILL19760x64220 (
);

FILL FILL_1__18190_ (
);

FILL FILL373920x217360 (
);

FILL FILL_1__9379_ (
);

FILL FILL_1__10697_ (
);

OR2X2 _9390_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_485_)
);

FILL FILL_0__15916_ (
);

FILL FILL262200x0 (
);

OR2X2 _18673_ (
    .A(_7578_),
    .B(_7575_),
    .Y(_7579_)
);

FILL FILL_0__18388_ (
);

OR2X2 _18253_ (
    .A(_7133_),
    .B(_7165_),
    .Y(_7166_)
);

FILL FILL358720x296400 (
);

FILL FILL249280x44460 (
);

FILL FILL476520x59280 (
);

FILL FILL_0__8489_ (
);

FILL FILL_0__9430_ (
);

FILL FILL_0__11836_ (
);

FILL FILL_0__9010_ (
);

OR2X2 _11701_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .B(_1718__bF$buf4),
    .Y(_1666_)
);

OR2X2 _19458_ (
    .A(gnd),
    .B(_8385__bF$buf0),
    .Y(_8341_)
);

OR2X2 _19038_ (
    .A(_7937_),
    .B(_7936_),
    .Y(_7938_)
);

AND2X2 _14593_ (
    .A(_3801_),
    .B(_3800_),
    .Y(_3738_[31])
);

OR2X2 _14173_ (
    .A(MemToReg_bF$buf4),
    .B(ALUOut[10]),
    .Y(_3560_)
);

OR2X2 _8908_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .B(_266__bF$buf2),
    .Y(_244_)
);

FILL FILL134520x247000 (
);

FILL FILL504640x326040 (
);

FILL FILL12920x247000 (
);

FILL FILL_1_BUFX2_insert360 (
);

FILL FILL18240x321100 (
);

NAND3X1 _12906_ (
    .A(_2266_),
    .B(\datapath_1.alu_1.ALUInA [22]),
    .C(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2471_)
);

FILL FILL_1_BUFX2_insert362 (
);

OR2X2 _15798_ (
    .A(_4744_),
    .B(_4747_),
    .Y(_4748_)
);

AND2X2 _15378_ (
    .A(_4223__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_4334_)
);

FILL FILL17480x88920 (
);

OR2X2 _10093_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .B(_860__bF$buf4),
    .Y(_854_)
);

FILL FILL_0__16874_ (
);

FILL FILL_0__16454_ (
);

FILL FILL196840x133380 (
);

FILL FILL177840x291460 (
);

OR2X2 _8661_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_119_)
);

FILL FILL323760x49400 (
);

FILL FILL221160x345800 (
);

FILL FILL_1__18666_ (
);

OR2X2 _11298_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_1457_)
);

FILL FILL_1__13381_ (
);

OR2X2 _17944_ (
    .A(_6860_),
    .B(_6857_),
    .Y(_6861_)
);

FILL FILL_0__17239_ (
);

OR2X2 _17524_ (
    .A(_6446_),
    .B(_6447_),
    .Y(_6448_)
);

OR2X2 _17104_ (
    .A(_6032_),
    .B(_6029_),
    .Y(_6033_)
);

FILL FILL_0__18600_ (
);

DFFSR _9866_ (
    .CLK(clk_bF$buf73),
    .D(_663_[23]),
    .Q(\datapath_1.regfile_1.regOut[11] [23]),
    .R(rst_bF$buf39),
    .S(vdd)
);

AND2X2 _9446_ (
    .A(_522_),
    .B(_521_),
    .Y(_465_[28])
);

AND2X2 _9026_ (
    .A(_302_),
    .B(_301_),
    .Y(_267_[17])
);

FILL FILL78280x281580 (
);

AND2X2 _18729_ (
    .A(_6236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_7634_)
);

FILL FILL245480x9880 (
);

AND2X2 _18309_ (
    .A(_6229__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_7221_)
);

FILL FILL_0__13999_ (
);

FILL FILL_0__13579_ (
);

OR2X2 _13864_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [16]),
    .Y(_3309_)
);

AND2X2 _13444_ (
    .A(_2976_),
    .B(_2975_),
    .Y(_2977_)
);

AOI21X1 _13024_ (
    .A(_2335_),
    .B(_2581_),
    .C(_2582_),
    .Y(_2583_)
);

FILL FILL78280x79040 (
);

FILL FILL_0__14940_ (
);

FILL FILL69160x256880 (
);

FILL FILL_0__9906_ (
);

FILL FILL_1__10086_ (
);

OR2X2 _14649_ (
    .A(\datapath_1.rd1 [7]),
    .B(_3869__bF$buf3),
    .Y(_3819_)
);

AND2X2 _14229_ (
    .A(_3597_),
    .B(_3596_),
    .Y(\datapath_1.mux_wd3.dout [28])
);

FILL FILL471960x14820 (
);

FILL FILL_1__16312_ (
);

FILL FILL_0__15305_ (
);

FILL FILL_0__10860_ (
);

FILL FILL_0__18197_ (
);

AND2X2 _18482_ (
    .A(_6293__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_7391_)
);

AND2X2 _18062_ (
    .A(_6289__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_6977_)
);

FILL FILL143640x365560 (
);

OR2X2 _10989_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_1311_)
);

FILL FILL_1__17517_ (
);

OR2X2 _10569_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_1091_)
);

OR2X2 _10149_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_871_)
);

DFFSR _11930_ (
    .CLK(clk_bF$buf25),
    .D(_1719_[23]),
    .Q(\datapath_1.regfile_1.regOut[27] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

AND2X2 _11510_ (
    .A(_1578_),
    .B(_1577_),
    .Y(_1521_[28])
);

FILL FILL_0__11225_ (
);

OR2X2 _19267_ (
    .A(_8163_),
    .B(_8162_),
    .Y(_8164_)
);

FILL FILL230280x276640 (
);

AND2X2 _8717_ (
    .A(_136_),
    .B(_199_),
    .Y(_135_[0])
);

FILL FILL367840x202540 (
);

FILL FILL471200x138320 (
);

AND2X2 _12715_ (
    .A(_2278_),
    .B(_2279_),
    .Y(_2280_)
);

FILL FILL479560x158080 (
);

FILL FILL198360x103740 (
);

FILL FILL_1_BUFX2_insert31 (
);

NAND2X1 _15187_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_4145_)
);

FILL FILL278920x365560 (
);

FILL FILL_1__17270_ (
);

FILL FILL_1_BUFX2_insert39 (
);

FILL FILL_1__8459_ (
);

FILL FILL_0__16263_ (
);

FILL FILL192280x256880 (
);

FILL FILL_1__9820_ (
);

FILL FILL275880x0 (
);

OR2X2 _8890_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .B(_266__bF$buf0),
    .Y(_232_)
);

OR2X2 _8470_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .B(_68__bF$buf2),
    .Y(_12_)
);

FILL FILL452960x88920 (
);

FILL FILL65360x286520 (
);

FILL FILL_0__17888_ (
);

FILL FILL388360x360620 (
);

FILL FILL_0__17468_ (
);

AND2X2 _17753_ (
    .A(_6300__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_6673_)
);

AND2X2 _17333_ (
    .A(_6258_),
    .B(_6219_),
    .Y(_6259_)
);

FILL FILL414200x355680 (
);

OR2X2 _9675_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_635_)
);

OR2X2 _9255_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_415_)
);

FILL FILL351120x103740 (
);

FILL FILL_0__8930_ (
);

FILL FILL_0__10916_ (
);

FILL FILL_0__8510_ (
);

FILL FILL93480x49400 (
);

OR2X2 _18958_ (
    .A(_7855_),
    .B(_7859_),
    .Y(_7860_)
);

AND2X2 _18538_ (
    .A(_6312__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_7446_)
);

AND2X2 _18118_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_7033_)
);

FILL FILL_1_BUFX2_insert1121 (
);

OR2X2 _13673_ (
    .A(_3156_),
    .B(_3155_),
    .Y(_3157_)
);

AOI21X1 _13253_ (
    .A(_2235_),
    .B(_2504_),
    .C(_2797_),
    .Y(_2798_)
);

FILL FILL428640x316160 (
);

FILL FILL_1_BUFX2_insert1129 (
);

FILL FILL329080x212420 (
);

FILL FILL42560x311220 (
);

FILL FILL352640x0 (
);

FILL FILL23560x148200 (
);

FILL FILL346560x222300 (
);

DFFSR _14878_ (
    .CLK(clk_bF$buf58),
    .D(_3870_[26]),
    .Q(_2_[26]),
    .R(rst_bF$buf104),
    .S(vdd)
);

AND2X2 _14458_ (
    .A(_3731_),
    .B(_3730_),
    .Y(_3672_[29])
);

AND2X2 _14038_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3452_)
);

FILL FILL_1__16961_ (
);

FILL FILL_0__15954_ (
);

FILL FILL_0__15534_ (
);

FILL FILL_0__15114_ (
);

FILL FILL177080x123500 (
);

AND2X2 _18291_ (
    .A(_6232__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_7203_)
);

FILL FILL110960x158080 (
);

OR2X2 _10798_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .B(_1256__bF$buf0),
    .Y(_1204_)
);

DFFSR _10378_ (
    .CLK(clk_bF$buf60),
    .D(_927_[19]),
    .Q(\datapath_1.regfile_1.regOut[15] [19]),
    .R(rst_bF$buf101),
    .S(vdd)
);

FILL FILL162640x345800 (
);

FILL FILL_0__16739_ (
);

OR2X2 _16604_ (
    .A(_5540_),
    .B(_5539_),
    .Y(_5541_)
);

FILL FILL_0__16319_ (
);

FILL FILL_0__11874_ (
);

FILL FILL76760x330980 (
);

OR2X2 _19496_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_8366_)
);

OR2X2 _19076_ (
    .A(_7974_),
    .B(_7975_),
    .Y(_7976_)
);

FILL FILL311600x330980 (
);

DFFSR _8946_ (
    .CLK(clk_bF$buf49),
    .D(_201_[6]),
    .Q(\datapath_1.regfile_1.regOut[4] [6]),
    .R(rst_bF$buf66),
    .S(vdd)
);

OR2X2 _8526_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_49_)
);

FILL FILL209000x9880 (
);

FILL FILL_1__13246_ (
);

AND2X2 _17809_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_6728_)
);

FILL FILL_1_BUFX2_insert741 (
);

XOR2X1 _12944_ (
    .A(_2167_),
    .B(_2489_),
    .Y(_2508_)
);

FILL FILL_0__12239_ (
);

NOR2X1 _12524_ (
    .A(_2113_),
    .B(\control_1.op [1]),
    .Y(_2114_)
);

AND2X2 _12104_ (
    .A(_1874_),
    .B(_1873_),
    .Y(_1851_[11])
);

FILL FILL498560x138320 (
);

FILL FILL15960x163020 (
);

FILL FILL234080x316160 (
);

FILL FILL_0__16492_ (
);

OR2X2 _13729_ (
    .A(_3204_),
    .B(_3203_),
    .Y(_3205_)
);

INVX1 _13309_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .Y(_2850_)
);

FILL FILL_1__15812_ (
);

FILL FILL_0__14805_ (
);

FILL FILL_1__18284_ (
);

BUFX2 BUFX2_insert410 (
    .A(_4172_),
    .Y(_4172__bF$buf0)
);

BUFX2 BUFX2_insert411 (
    .A(_4228_),
    .Y(_4228__bF$buf4)
);

BUFX2 BUFX2_insert412 (
    .A(_4228_),
    .Y(_4228__bF$buf3)
);

BUFX2 BUFX2_insert413 (
    .A(_4228_),
    .Y(_4228__bF$buf2)
);

OR2X2 _17982_ (
    .A(_6898_),
    .B(_6897_),
    .Y(_6899_)
);

BUFX2 BUFX2_insert414 (
    .A(_4228_),
    .Y(_4228__bF$buf1)
);

AND2X2 _17562_ (
    .A(_6262__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_6485_)
);

BUFX2 BUFX2_insert415 (
    .A(_4228_),
    .Y(_4228__bF$buf0)
);

FILL FILL_0__17277_ (
);

BUFX2 BUFX2_insert416 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf4 )
);

OR2X2 _17142_ (
    .A(_6070_),
    .B(_6067_),
    .Y(_6071_)
);

BUFX2 BUFX2_insert417 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf3 )
);

BUFX2 BUFX2_insert418 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf2 )
);

BUFX2 BUFX2_insert419 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf1 )
);

FILL FILL51680x108680 (
);

DFFSR _9484_ (
    .CLK(clk_bF$buf74),
    .D(_465_[28]),
    .Q(\datapath_1.regfile_1.regOut[8] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

OR2X2 _9064_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .B(_332__bF$buf2),
    .Y(_328_)
);

FILL FILL433200x335920 (
);

FILL FILL_1__19489_ (
);

FILL FILL19760x271700 (
);

FILL FILL_0__10305_ (
);

AND2X2 _18767_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_7672_)
);

OR2X2 _18347_ (
    .A(_7256_),
    .B(_7257_),
    .Y(_7258_)
);

FILL FILL_0__13197_ (
);

OR2X2 _13482_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [21]),
    .Y(_3011_)
);

AND2X2 _13062_ (
    .A(_2618_),
    .B(_2263_),
    .Y(_2619_)
);

FILL FILL336680x177840 (
);

FILL FILL_0__19423_ (
);

FILL FILL_0__19003_ (
);

FILL FILL_1__12517_ (
);

FILL FILL_0__9944_ (
);

FILL FILL_0__9104_ (
);

OR2X2 _14687_ (
    .A(vdd),
    .B(\datapath_1.a [20]),
    .Y(_3844_)
);

OR2X2 _14267_ (
    .A(vdd),
    .B(ALUOut[9]),
    .Y(_3624_)
);

FILL FILL490960x247000 (
);

FILL FILL_0__15763_ (
);

FILL FILL_0__15343_ (
);

FILL FILL421800x108680 (
);

FILL FILL112480x128440 (
);

FILL FILL152000x237120 (
);

FILL FILL_1__8900_ (
);

FILL FILL186960x59280 (
);

AND2X2 _10187_ (
    .A(_896_),
    .B(_895_),
    .Y(_861_[17])
);

FILL FILL_1__17135_ (
);

FILL FILL_1__12270_ (
);

FILL FILL_0__16968_ (
);

OR2X2 _16833_ (
    .A(_5765_),
    .B(_5762_),
    .Y(_5766_)
);

AND2X2 _16413_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_5353_)
);

FILL FILL_0__11683_ (
);

FILL FILL233320x167960 (
);

OR2X2 _8755_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .B(_200__bF$buf1),
    .Y(_162_)
);

FILL FILL451440x291460 (
);

FILL FILL38000x355680 (
);

FILL FILL503880x138320 (
);

FILL FILL_1__13895_ (
);

FILL FILL_1__13475_ (
);

AND2X2 _17618_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_6540_)
);

NOR2X1 _12753_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2318_)
);

FILL FILL_0__12468_ (
);

OR2X2 _12333_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_1987_)
);

FILL FILL201400x301340 (
);

FILL FILL370880x212420 (
);

OR2X2 _13958_ (
    .A(_3383_),
    .B(_3382_),
    .Y(_3384_)
);

FILL FILL351880x370500 (
);

OR2X2 _13538_ (
    .A(ALUOut[16]),
    .B(_3079__bF$buf2),
    .Y(_3047_)
);

OR2X2 _13118_ (
    .A(_2157__bF$buf2),
    .B(_2670_),
    .Y(_2671_)
);

FILL FILL281960x375440 (
);

OR2X2 _17791_ (
    .A(_6710_),
    .B(_6709_),
    .Y(_6711_)
);

AND2X2 _17371_ (
    .A(_6296_),
    .B(_6209_),
    .Y(_6297_)
);

FILL FILL_0__17086_ (
);

FILL FILL505400x306280 (
);

AND2X2 _9293_ (
    .A(_440_),
    .B(_439_),
    .Y(_399_[20])
);

FILL FILL_1__11961_ (
);

FILL FILL_0__15819_ (
);

OR2X2 _18996_ (
    .A(_7896_),
    .B(_7895_),
    .Y(_7897_)
);

OR2X2 _18576_ (
    .A(_7483_),
    .B(_7476_),
    .Y(_7484_)
);

AND2X2 _18156_ (
    .A(_6259__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_7070_)
);

FILL FILL422560x54340 (
);

AND2X2 _13291_ (
    .A(_2833_),
    .B(_2828_),
    .Y(_2834_)
);

FILL FILL130720x83980 (
);

FILL FILL82080x59280 (
);

FILL FILL215080x54340 (
);

FILL FILL_1__12326_ (
);

FILL FILL161120x355680 (
);

FILL FILL_0__9753_ (
);

FILL FILL_0__11739_ (
);

FILL FILL_0__11319_ (
);

OR2X2 _11604_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_1621_)
);

DFFSR _14496_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[31]),
    .Q(\datapath_1.Data [31]),
    .R(rst_bF$buf85),
    .S(vdd)
);

AND2X2 _14076_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3485_)
);

FILL FILL49400x123500 (
);

FILL FILL_0__15992_ (
);

FILL FILL_0__15572_ (
);

NAND2X1 _12809_ (
    .A(ALUControl[2]),
    .B(_2155_),
    .Y(_2374_)
);

FILL FILL42560x14820 (
);

FILL FILL_1__17784_ (
);

AND2X2 _16642_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_5578_)
);

FILL FILL_0__16357_ (
);

AND2X2 _16222_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_5165_)
);

FILL FILL_0__11492_ (
);

AND2X2 _8984_ (
    .A(_274_),
    .B(_273_),
    .Y(_267_[3])
);

DFFSR _8564_ (
    .CLK(clk_bF$buf45),
    .D(_3_[11]),
    .Q(\datapath_1.regfile_1.regOut[1] [11]),
    .R(rst_bF$buf54),
    .S(vdd)
);

AND2X2 _17847_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_6766_)
);

AND2X2 _17427_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_6352_)
);

FILL FILL315400x321100 (
);

FILL FILL69920x14820 (
);

OR2X2 _17007_ (
    .A(_5934_),
    .B(_5937_),
    .Y(_5938_)
);

FILL FILL_0__12697_ (
);

OR2X2 _12982_ (
    .A(_2540_),
    .B(_2542_),
    .Y(_2543_)
);

FILL FILL_0__12277_ (
);

AND2X2 _12562_ (
    .A(_2082_),
    .B(_2081_),
    .Y(_2083_)
);

OR2X2 _12142_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .B(_1916__bF$buf4),
    .Y(_1900_)
);

FILL FILL_0__18923_ (
);

FILL FILL_0__18503_ (
);

OR2X2 _9769_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .B(_728__bF$buf1),
    .Y(_678_)
);

FILL FILL47880x74100 (
);

DFFSR _9349_ (
    .CLK(clk_bF$buf72),
    .D(_399_[22]),
    .Q(\datapath_1.regfile_1.regOut[7] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

AND2X2 _13767_ (
    .A(_3084__bF$buf2),
    .B(\datapath_1.PCJump [25]),
    .Y(_3237_)
);

NAND3X1 _13347_ (
    .A(_2886_),
    .B(_2547_),
    .C(_2874_),
    .Y(_2887_)
);

FILL FILL_1__15430_ (
);

FILL FILL_0__14423_ (
);

FILL FILL_0__14003_ (
);

OR2X2 _17180_ (
    .A(_6107_),
    .B(_6106_),
    .Y(_6108_)
);

FILL FILL432440x330980 (
);

FILL FILL_1__16635_ (
);

FILL FILL253840x24700 (
);

FILL FILL_0__15628_ (
);

AND2X2 _15913_ (
    .A(_4241__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_4861_)
);

FILL FILL_0__15208_ (
);

FILL FILL80560x79040 (
);

FILL FILL294120x217360 (
);

FILL FILL323000x54340 (
);

AND2X2 _18385_ (
    .A(_7295_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd1 [15])
);

FILL FILL467400x237120 (
);

FILL FILL_0__19041_ (
);

FILL FILL180120x335920 (
);

FILL FILL_0__11968_ (
);

FILL FILL_0__9562_ (
);

FILL FILL_0__9142_ (
);

OR2X2 _11833_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .B(_1784__bF$buf1),
    .Y(_1734_)
);

DFFSR _11413_ (
    .CLK(clk_bF$buf74),
    .D(_1455_[22]),
    .Q(\datapath_1.regfile_1.regOut[23] [22]),
    .R(rst_bF$buf47),
    .S(vdd)
);

FILL FILL_0__11128_ (
);

FILL FILL_0__15381_ (
);

FILL FILL256880x197600 (
);

OR2X2 _12618_ (
    .A(_2182_),
    .B(_2172_),
    .Y(_2183_)
);

FILL FILL_1__14701_ (
);

FILL FILL_0__16586_ (
);

OR2X2 _16871_ (
    .A(_5803_),
    .B(_5800_),
    .Y(_5804_)
);

AND2X2 _16451_ (
    .A(_4210__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_5390_)
);

OR2X2 _16031_ (
    .A(_4976_),
    .B(_4975_),
    .Y(_4977_)
);

FILL FILL305520x276640 (
);

FILL FILL50920x163020 (
);

OR2X2 _8793_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_187_)
);

FILL FILL381520x54340 (
);

FILL FILL146680x217360 (
);

AND2X2 _17656_ (
    .A(_6216__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_6578_)
);

AND2X2 _17236_ (
    .A(_4181__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_6163_)
);

NOR2X1 _12791_ (
    .A(_2355_),
    .B(_2353_),
    .Y(_2356_)
);

AND2X2 _12371_ (
    .A(_2012_),
    .B(_2011_),
    .Y(_1983_[14])
);

FILL FILL_0__12086_ (
);

FILL FILL_0__18732_ (
);

DFFSR _9998_ (
    .CLK(clk_bF$buf55),
    .D(_729_[26]),
    .Q(\datapath_1.regfile_1.regOut[12] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

AND2X2 _9578_ (
    .A(_590_),
    .B(_589_),
    .Y(_531_[29])
);

AND2X2 _9158_ (
    .A(_370_),
    .B(_369_),
    .Y(_333_[18])
);

FILL FILL56240x103740 (
);

FILL FILL_0__10819_ (
);

FILL FILL_0_BUFX2_insert780 (
);

FILL FILL_0_BUFX2_insert781 (
);

FILL FILL_0_BUFX2_insert782 (
);

FILL FILL_0_BUFX2_insert783 (
);

AND2X2 _13996_ (
    .A(_3347__bF$buf1),
    .B(\datapath_1.PCJump [13]),
    .Y(_3416_)
);

FILL FILL_0_BUFX2_insert784 (
);

OR2X2 _13576_ (
    .A(IorD_bF$buf0),
    .B(\datapath_1.PCJump [29]),
    .Y(_3072_)
);

OAI21X1 _13156_ (
    .A(_2210_),
    .B(_2225_),
    .C(_2258_),
    .Y(_2707_)
);

FILL FILL_0_BUFX2_insert786 (
);

FILL FILL_0_BUFX2_insert788 (
);

FILL FILL_0__19517_ (
);

FILL FILL_0__14652_ (
);

FILL FILL_0__14232_ (
);

FILL FILL_0__15857_ (
);

FILL FILL_0__15437_ (
);

AND2X2 _15722_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_4673_)
);

AND2X2 _15302_ (
    .A(_4217__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_4259_)
);

FILL FILL_0__10992_ (
);

FILL FILL_0__10572_ (
);

FILL FILL71440x187720 (
);

AND2X2 _18194_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_7107_)
);

FILL FILL_0__19270_ (
);

FILL FILL_1__17649_ (
);

OR2X2 _16927_ (
    .A(_5857_),
    .B(_5858_),
    .Y(_5859_)
);

AND2X2 _16507_ (
    .A(_4236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_5445_)
);

FILL FILL_0__9791_ (
);

FILL FILL_0__9371_ (
);

AND2X2 _11642_ (
    .A(_1646_),
    .B(_1645_),
    .Y(_1587_[29])
);

AND2X2 _11222_ (
    .A(_1426_),
    .B(_1425_),
    .Y(_1389_[18])
);

AND2X2 _19399_ (
    .A(_6302__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_8294_)
);

AND2X2 _8849_ (
    .A(_204_),
    .B(_203_),
    .Y(_201_[1])
);

BUFX2 _8429_ (
    .A(_2_[5]),
    .Y(memoryWriteData[5])
);

FILL FILL_1__13989_ (
);

FILL FILL329080x59280 (
);

FILL FILL142880x247000 (
);

FILL FILL346560x182780 (
);

NAND3X1 _12847_ (
    .A(_2411_),
    .B(\datapath_1.alu_1.ALUInB [6]),
    .C(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2412_)
);

DFFSR _12427_ (
    .CLK(clk_bF$buf79),
    .D(_1983_[4]),
    .Q(\datapath_1.regfile_1.regOut[31] [4]),
    .R(rst_bF$buf2),
    .S(vdd)
);

OR2X2 _12007_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .B(_1850__bF$buf4),
    .Y(_1830_)
);

FILL FILL_1__14510_ (
);

FILL FILL_0__13923_ (
);

FILL FILL_0__13503_ (
);

FILL FILL282720x128440 (
);

FILL FILL_0__16395_ (
);

OR2X2 _16680_ (
    .A(_5608_),
    .B(_5615_),
    .Y(_5616_)
);

OR2X2 _16260_ (
    .A(_5201_),
    .B(_5200_),
    .Y(_5202_)
);

FILL FILL_1__9952_ (
);

FILL FILL_1__10850_ (
);

FILL FILL117800x69160 (
);

FILL FILL_0__14708_ (
);

OR2X2 _17885_ (
    .A(_6802_),
    .B(_6801_),
    .Y(_6803_)
);

FILL FILL103360x291460 (
);

AND2X2 _17465_ (
    .A(_6326__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_6390_)
);

AND2X2 _17045_ (
    .A(_4135__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_5975_)
);

DFFSR _12180_ (
    .CLK(clk_bF$buf39),
    .D(_1851_[15]),
    .Q(\datapath_1.regfile_1.regOut[29] [15]),
    .R(rst_bF$buf69),
    .S(vdd)
);

FILL FILL360240x335920 (
);

FILL FILL_0__18121_ (
);

OR2X2 _9387_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_483_)
);

FILL FILL_1__11215_ (
);

FILL FILL_0__8642_ (
);

AND2X2 _10913_ (
    .A(_1260_),
    .B(_1259_),
    .Y(_1257_[1])
);

FILL FILL_0__10208_ (
);

FILL FILL199880x350740 (
);

FILL FILL231040x326040 (
);

OR2X2 _13385_ (
    .A(_2157__bF$buf1),
    .B(_2921_),
    .Y(_2922_)
);

FILL FILL293360x0 (
);

FILL FILL193040x24700 (
);

FILL FILL413440x237120 (
);

FILL FILL322240x19760 (
);

FILL FILL_0__9007_ (
);

FILL FILL_1__16253_ (
);

FILL FILL174800x237120 (
);

OR2X2 _15951_ (
    .A(_4897_),
    .B(_4896_),
    .Y(_4898_)
);

OR2X2 _15531_ (
    .A(_4484_),
    .B(_4483_),
    .Y(_4485_)
);

AND2X2 _15111_ (
    .A(_4090_),
    .B(_4084_),
    .Y(_4091_)
);

FILL FILL280440x311220 (
);

FILL FILL193800x98800 (
);

FILL FILL_1__8803_ (
);

FILL FILL_1__12593_ (
);

FILL FILL278160x291460 (
);

OR2X2 _16736_ (
    .A(_5667_),
    .B(_5670_),
    .Y(_5671_)
);

AND2X2 _16316_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_5257_)
);

OR2X2 _11871_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_1759_)
);

FILL FILL_0__9180_ (
);

OR2X2 _11451_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_1539_)
);

FILL FILL_0__11166_ (
);

DFFSR _11031_ (
    .CLK(clk_bF$buf104),
    .D(_1257_[27]),
    .Q(\datapath_1.regfile_1.regOut[20] [27]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL447640x256880 (
);

FILL FILL370120x0 (
);

FILL FILL327560x79040 (
);

OR2X2 _8658_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_117_)
);

FILL FILL61560x251940 (
);

FILL FILL92720x237120 (
);

XNOR2X1 _12656_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2221_)
);

AND2X2 _12236_ (
    .A(_1942_),
    .B(_1941_),
    .Y(_1917_[12])
);

FILL FILL197600x98800 (
);

FILL FILL_0__13732_ (
);

FILL FILL_0__13312_ (
);

FILL FILL295640x167960 (
);

FILL FILL_0_BUFX2_insert1131 (
);

FILL FILL_0_BUFX2_insert1133 (
);

FILL FILL_0_BUFX2_insert1135 (
);

FILL FILL_0_BUFX2_insert1136 (
);

FILL FILL_0_BUFX2_insert1137 (
);

FILL FILL_0_BUFX2_insert1138 (
);

FILL FILL_1__9761_ (
);

FILL FILL_0_BUFX2_insert1139 (
);

FILL FILL_1__15104_ (
);

FILL FILL166440x158080 (
);

FILL FILL_0__14937_ (
);

OR2X2 _14802_ (
    .A(\datapath_1.rd2 [15]),
    .B(_3935__bF$buf2),
    .Y(_3901_)
);

FILL FILL_0__14517_ (
);

FILL FILL348080x29640 (
);

OR2X2 _17694_ (
    .A(_6614_),
    .B(_6613_),
    .Y(_6615_)
);

AND2X2 _17274_ (
    .A(_6200_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [31])
);

FILL FILL152760x182780 (
);

FILL FILL_0__18770_ (
);

FILL FILL_0__18350_ (
);

FILL FILL_1__16729_ (
);

OR2X2 _9196_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .B(_398__bF$buf1),
    .Y(_396_)
);

FILL FILL_0__8871_ (
);

FILL FILL_0__8451_ (
);

FILL FILL_0__10857_ (
);

FILL FILL259160x103740 (
);

FILL FILL_0__10437_ (
);

OR2X2 _10722_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_1173_)
);

FILL FILL_0__10017_ (
);

OR2X2 _10302_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_953_)
);

OR2X2 _18899_ (
    .A(_7800_),
    .B(_7801_),
    .Y(_7802_)
);

OR2X2 _18479_ (
    .A(_7387_),
    .B(_7380_),
    .Y(_7388_)
);

OR2X2 _18059_ (
    .A(_6940_),
    .B(_6974_),
    .Y(_6975_)
);

OR2X2 _13194_ (
    .A(_2428_),
    .B(_2415_),
    .Y(_2743_)
);

FILL FILL204440x64220 (
);

FILL FILL221160x14820 (
);

FILL FILL58520x217360 (
);

FILL FILL_0__19555_ (
);

OR2X2 _19420_ (
    .A(_8311_),
    .B(_8314_),
    .Y(_8315_)
);

FILL FILL_0__19135_ (
);

FILL FILL6080x158080 (
);

AND2X2 _19000_ (
    .A(_6282__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [25]),
    .Y(_7901_)
);

FILL FILL471200x251940 (
);

DFFSR _11927_ (
    .CLK(clk_bF$buf56),
    .D(_1719_[20]),
    .Q(\datapath_1.regfile_1.regOut[27] [20]),
    .R(rst_bF$buf49),
    .S(vdd)
);

AND2X2 _11507_ (
    .A(_1576_),
    .B(_1575_),
    .Y(_1521_[27])
);

FILL FILL205200x182780 (
);

OR2X2 _14399_ (
    .A(vdd),
    .B(\datapath_1.Data [10]),
    .Y(_3692_)
);

FILL FILL449160x360620 (
);

FILL FILL115520x316160 (
);

FILL FILL_0__15475_ (
);

OR2X2 _15760_ (
    .A(_4706_),
    .B(_4709_),
    .Y(_4710_)
);

FILL FILL_0__15055_ (
);

AND2X2 _15340_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_4297_)
);

FILL FILL_0__10190_ (
);

FILL FILL101840x340860 (
);

AND2X2 _16965_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_5896_)
);

AND2X2 _16545_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_5483_)
);

OR2X2 _16125_ (
    .A(_5067_),
    .B(_5068_),
    .Y(_5069_)
);

DFFSR _11680_ (
    .CLK(clk_bF$buf27),
    .D(_1587_[31]),
    .Q(\datapath_1.regfile_1.regOut[25] [31]),
    .R(rst_bF$buf28),
    .S(vdd)
);

FILL FILL342000x108680 (
);

OR2X2 _11260_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .B(_1454__bF$buf3),
    .Y(_1452_)
);

FILL FILL_0__17621_ (
);

FILL FILL_0__17201_ (
);

FILL FILL135280x49400 (
);

OR2X2 _8887_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .B(_266__bF$buf2),
    .Y(_230_)
);

OR2X2 _8467_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .B(_68__bF$buf0),
    .Y(_10_)
);

FILL FILL33440x316160 (
);

NAND3X1 _12885_ (
    .A(_2262_),
    .B(_2263_),
    .C(_2267_),
    .Y(_2450_)
);

FILL FILL_1__19413_ (
);

AND2X2 _12465_ (
    .A(_2049_),
    .B(\aluControl_1.inst [2]),
    .Y(_2058_)
);

DFFSR _12045_ (
    .CLK(clk_bF$buf24),
    .D(_1785_[9]),
    .Q(\datapath_1.regfile_1.regOut[28] [9]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_0__13961_ (
);

FILL FILL_0__13121_ (
);

FILL FILL262960x281580 (
);

FILL FILL443080x301340 (
);

FILL FILL_1_BUFX2_insert3 (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_0__8927_ (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1__9570_ (
);

FILL FILL346560x49400 (
);

FILL FILL_1_BUFX2_insert1093 (
);

FILL FILL223440x345800 (
);

FILL FILL253840x256880 (
);

FILL FILL_1_BUFX2_insert1095 (
);

FILL FILL_1_BUFX2_insert1097 (
);

FILL FILL_1__15753_ (
);

FILL FILL_0__14326_ (
);

DFFSR _14611_ (
    .CLK(clk_bF$buf65),
    .D(_3738_[17]),
    .Q(\datapath_1.PCJump [19]),
    .R(rst_bF$buf91),
    .S(vdd)
);

AND2X2 _17083_ (
    .A(_4195__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_6012_)
);

FILL FILL376200x44460 (
);

FILL FILL_1__16118_ (
);

OR2X2 _15816_ (
    .A(_4764_),
    .B(_4761_),
    .Y(_4765_)
);

FILL FILL_0__8680_ (
);

OR2X2 _10951_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .B(_1322__bF$buf0),
    .Y(_1286_)
);

FILL FILL_0__10666_ (
);

OR2X2 _10531_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .B(_1124__bF$buf4),
    .Y(_1066_)
);

DFFSR _10111_ (
    .CLK(clk_bF$buf88),
    .D(_795_[10]),
    .Q(\datapath_1.regfile_1.regOut[13] [10]),
    .R(rst_bF$buf95),
    .S(vdd)
);

AND2X2 _18288_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_7200_)
);

FILL FILL_0__19364_ (
);

FILL FILL_1__12878_ (
);

FILL FILL_1__12458_ (
);

FILL FILL_0__9885_ (
);

OR2X2 _11736_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_1689_)
);

FILL FILL_0__9045_ (
);

OR2X2 _11316_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_1469_)
);

FILL FILL436240x4940 (
);

FILL FILL435480x98800 (
);

FILL FILL145920x365560 (
);

FILL FILL_1__17076_ (
);

FILL FILL471960x88920 (
);

AND2X2 _16774_ (
    .A(_4217__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_5708_)
);

FILL FILL232560x276640 (
);

FILL FILL_0__16069_ (
);

AND2X2 _16354_ (
    .A(_4146__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_5295_)
);

FILL FILL_0__17850_ (
);

FILL FILL264480x88920 (
);

FILL FILL_0__17010_ (
);

DFFSR _8696_ (
    .CLK(clk_bF$buf63),
    .D(_69_[14]),
    .Q(\datapath_1.regfile_1.regOut[2] [14]),
    .R(rst_bF$buf4),
    .S(vdd)
);

BUFX2 BUFX2_insert380 (
    .A(_6262_),
    .Y(_6262__bF$buf0)
);

BUFX2 BUFX2_insert381 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf4 )
);

BUFX2 BUFX2_insert382 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf3 )
);

BUFX2 BUFX2_insert383 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf2 )
);

OR2X2 _17979_ (
    .A(_6894_),
    .B(_6895_),
    .Y(_6896_)
);

BUFX2 BUFX2_insert384 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf1 )
);

BUFX2 BUFX2_insert385 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf0 )
);

OR2X2 _17559_ (
    .A(_6480_),
    .B(_6481_),
    .Y(_6482_)
);

BUFX2 BUFX2_insert386 (
    .A(_6259_),
    .Y(_6259__bF$buf4)
);

AND2X2 _17139_ (
    .A(_4158__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_6068_)
);

BUFX2 BUFX2_insert387 (
    .A(_6259_),
    .Y(_6259__bF$buf3)
);

BUFX2 BUFX2_insert388 (
    .A(_6259_),
    .Y(_6259__bF$buf2)
);

BUFX2 BUFX2_insert389 (
    .A(_6259_),
    .Y(_6259__bF$buf1)
);

AND2X2 _12694_ (
    .A(_2226_),
    .B(_2258_),
    .Y(_2259_)
);

OR2X2 _12274_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .B(_1982__bF$buf0),
    .Y(_1968_)
);

FILL FILL338200x74100 (
);

FILL FILL437760x271700 (
);

FILL FILL_0__18635_ (
);

OR2X2 _18920_ (
    .A(_7814_),
    .B(_7821_),
    .Y(_7822_)
);

FILL FILL_0__18215_ (
);

AND2X2 _18500_ (
    .A(_6255__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_7409_)
);

FILL FILL_0__13350_ (
);

FILL FILL_1__11309_ (
);

FILL FILL367840x276640 (
);

FILL FILL_0__8736_ (
);

FILL FILL126920x311220 (
);

AND2X2 _13899_ (
    .A(_3332_),
    .B(_3331_),
    .Y(\datapath_1.alu_1.ALUInA [27])
);

OR2X2 _13479_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [20]),
    .Y(_3009_)
);

OR2X2 _13059_ (
    .A(_2451_),
    .B(_2615_),
    .Y(_2616_)
);

FILL FILL_1__15982_ (
);

FILL FILL454480x187720 (
);

OR2X2 _14840_ (
    .A(vdd),
    .B(_2_[28]),
    .Y(_3926_)
);

FILL FILL_0__14555_ (
);

OR2X2 _14420_ (
    .A(vdd),
    .B(\datapath_1.Data [17]),
    .Y(_3706_)
);

OR2X2 _14000_ (
    .A(_3419_),
    .B(_3418_),
    .Y(_3420_)
);

FILL FILL213560x222300 (
);

FILL FILL448400x143260 (
);

FILL FILL308560x128440 (
);

FILL FILL353400x103740 (
);

FILL FILL_1__16767_ (
);

OR2X2 _15625_ (
    .A(_4569_),
    .B(_4576_),
    .Y(_4577_)
);

OR2X2 _15205_ (
    .A(_4162_),
    .B(_4156_),
    .Y(_4163_)
);

DFFSR _10760_ (
    .CLK(clk_bF$buf37),
    .D(_1125_[14]),
    .Q(\datapath_1.regfile_1.regOut[18] [14]),
    .R(rst_bF$buf103),
    .S(vdd)
);

AND2X2 _10340_ (
    .A(_978_),
    .B(_977_),
    .Y(_927_[25])
);

FILL FILL_0__10055_ (
);

FILL FILL334400x261820 (
);

OR2X2 _18097_ (
    .A(_7011_),
    .B(_7010_),
    .Y(_7012_)
);

FILL FILL_0__16701_ (
);

FILL FILL211280x296400 (
);

FILL FILL_0__19173_ (
);

FILL FILL25840x148200 (
);

FILL FILL348840x222300 (
);

FILL FILL361760x217360 (
);

FILL FILL44080x217360 (
);

FILL FILL_0__9694_ (
);

OR2X2 _11965_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .B(_1850__bF$buf4),
    .Y(_1802_)
);

FILL FILL_0__9274_ (
);

FILL FILL_1__18913_ (
);

DFFSR _11545_ (
    .CLK(clk_bF$buf16),
    .D(_1521_[25]),
    .Q(\datapath_1.regfile_1.regOut[24] [25]),
    .R(rst_bF$buf76),
    .S(vdd)
);

OR2X2 _11125_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .B(_1388__bF$buf1),
    .Y(_1382_)
);

FILL FILL_0__12621_ (
);

FILL FILL_0__12201_ (
);

FILL FILL120080x59280 (
);

FILL FILL_0__15093_ (
);

FILL FILL_1__8650_ (
);

FILL FILL_1__14413_ (
);

FILL FILL_0__13826_ (
);

FILL FILL457520x9880 (
);

OR2X2 _16583_ (
    .A(_5518_),
    .B(_5519_),
    .Y(_5520_)
);

FILL FILL_0__16298_ (
);

OR2X2 _16163_ (
    .A(_5105_),
    .B(_5106_),
    .Y(_5107_)
);

FILL FILL414200x217360 (
);

FILL FILL221920x9880 (
);

FILL FILL_1__15618_ (
);

OR2X2 _17788_ (
    .A(_6707_),
    .B(_6704_),
    .Y(_6708_)
);

AND2X2 _17368_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_6294_)
);

AND2X2 _12083_ (
    .A(_1860_),
    .B(_1859_),
    .Y(_1851_[4])
);

FILL FILL_1__19031_ (
);

FILL FILL236360x316160 (
);

FILL FILL323760x321100 (
);

FILL FILL_0__18864_ (
);

FILL FILL_0__18444_ (
);

FILL FILL_0__18024_ (
);

FILL FILL_0__8545_ (
);

OR2X2 _10816_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_1256__bF$buf4),
    .Y(_1216_)
);

FILL FILL107920x14820 (
);

FILL FILL495520x9880 (
);

AND2X2 _13288_ (
    .A(_2524_),
    .B(_2232_),
    .Y(_2831_)
);

FILL FILL_1__15371_ (
);

FILL FILL_0__19229_ (
);

OR2X2 _19514_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_8378_)
);

FILL FILL_0__14784_ (
);

FILL FILL226480x261820 (
);

FILL FILL467400x123500 (
);

FILL FILL363280x321100 (
);

FILL FILL231800x44460 (
);

FILL FILL_0__15989_ (
);

OR2X2 _15854_ (
    .A(_4801_),
    .B(_4802_),
    .Y(_4803_)
);

FILL FILL_0__15569_ (
);

FILL FILL_0__15149_ (
);

AND2X2 _15434_ (
    .A(_4189__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_4389_)
);

NAND2X1 _15014_ (
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_4003_)
);

FILL FILL_0__16510_ (
);

FILL FILL484120x360620 (
);

FILL FILL100320x167960 (
);

FILL FILL_1__12076_ (
);

AND2X2 _16639_ (
    .A(_4135__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_5575_)
);

AND2X2 _16219_ (
    .A(_4183__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_5162_)
);

AND2X2 _11774_ (
    .A(_1714_),
    .B(_1713_),
    .Y(_1653_[30])
);

AND2X2 _11354_ (
    .A(_1494_),
    .B(_1493_),
    .Y(_1455_[19])
);

FILL FILL_0__11069_ (
);

FILL FILL_0__17715_ (
);

FILL FILL_0__12850_ (
);

FILL FILL114760x128440 (
);

FILL FILL_0__12010_ (
);

OR2X2 _9922_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .B(_794__bF$buf4),
    .Y(_760_)
);

OR2X2 _9502_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_596__bF$buf1),
    .Y(_540_)
);

INVX1 _12979_ (
    .A(_2321_),
    .Y(_2540_)
);

INVX1 _12559_ (
    .A(_2111_),
    .Y(_2080_)
);

OR2X2 _12139_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_1916__bF$buf0),
    .Y(_1898_)
);

FILL FILL_1__14222_ (
);

AND2X2 _13920_ (
    .A(_3350__bF$buf1),
    .B(_2_[0]),
    .Y(_3351_)
);

FILL FILL_0__13215_ (
);

AND2X2 _13500_ (
    .A(_3021_),
    .B(_3020_),
    .Y(_1_[3])
);

FILL FILL235600x167960 (
);

FILL FILL162640x29640 (
);

OR2X2 _16392_ (
    .A(_5331_),
    .B(_5328_),
    .Y(_5332_)
);

FILL FILL_1__9664_ (
);

FILL FILL_1__15847_ (
);

FILL FILL_1__10982_ (
);

FILL FILL41040x251940 (
);

FILL FILL294880x232180 (
);

OR2X2 _14705_ (
    .A(vdd),
    .B(\datapath_1.a [26]),
    .Y(_3856_)
);

BUFX2 BUFX2_insert760 (
    .A(_1652_),
    .Y(_1652__bF$buf2)
);

FILL FILL444600x266760 (
);

BUFX2 BUFX2_insert761 (
    .A(_1652_),
    .Y(_1652__bF$buf1)
);

BUFX2 BUFX2_insert762 (
    .A(_1652_),
    .Y(_1652__bF$buf0)
);

BUFX2 BUFX2_insert763 (
    .A(_6326_),
    .Y(_6326__bF$buf4)
);

BUFX2 BUFX2_insert764 (
    .A(_6326_),
    .Y(_6326__bF$buf3)
);

FILL FILL212040x232180 (
);

AND2X2 _17597_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_6520_)
);

BUFX2 BUFX2_insert765 (
    .A(_6326_),
    .Y(_6326__bF$buf2)
);

BUFX2 BUFX2_insert766 (
    .A(_6326_),
    .Y(_6326__bF$buf1)
);

OR2X2 _17177_ (
    .A(_6089_),
    .B(_6104_),
    .Y(_6105_)
);

BUFX2 BUFX2_insert767 (
    .A(_6326_),
    .Y(_6326__bF$buf0)
);

BUFX2 BUFX2_insert768 (
    .A(_6229_),
    .Y(_6229__bF$buf4)
);

BUFX2 BUFX2_insert769 (
    .A(_6229_),
    .Y(_6229__bF$buf3)
);

FILL FILL249280x355680 (
);

FILL FILL_0__18673_ (
);

DFFSR _9099_ (
    .CLK(clk_bF$buf108),
    .D(_267_[30]),
    .Q(\datapath_1.regfile_1.regOut[5] [30]),
    .R(rst_bF$buf66),
    .S(vdd)
);

FILL FILL_1__11347_ (
);

FILL FILL_0__8774_ (
);

DFFSR _10625_ (
    .CLK(clk_bF$buf22),
    .D(_1059_[8]),
    .Q(\datapath_1.regfile_1.regOut[17] [8]),
    .R(rst_bF$buf74),
    .S(vdd)
);

AND2X2 _10205_ (
    .A(_908_),
    .B(_907_),
    .Y(_861_[23])
);

AND2X2 _13097_ (
    .A(_2651_),
    .B(_2646_),
    .Y(_2652_)
);

FILL FILL_0__11701_ (
);

FILL FILL_0__19458_ (
);

FILL FILL_0__19038_ (
);

OR2X2 _19323_ (
    .A(_8218_),
    .B(_8215_),
    .Y(_8219_)
);

FILL FILL_0__14173_ (
);

FILL FILL_0__9139_ (
);

FILL FILL370880x286520 (
);

FILL FILL_0__12906_ (
);

FILL FILL_0__15798_ (
);

FILL FILL421800x24700 (
);

FILL FILL_0__15378_ (
);

OR2X2 _15663_ (
    .A(_4611_),
    .B(_4614_),
    .Y(_4615_)
);

AND2X2 _15243_ (
    .A(_4200__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [0]),
    .Y(_4201_)
);

FILL FILL_1__8935_ (
);

FILL FILL247760x311220 (
);

AND2X2 _16868_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_5801_)
);

OR2X2 _16448_ (
    .A(_5385_),
    .B(_5386_),
    .Y(_5387_)
);

FILL FILL297920x44460 (
);

OR2X2 _16028_ (
    .A(_4973_),
    .B(_4972_),
    .Y(_4974_)
);

FILL FILL_1__18531_ (
);

FILL FILL_0__11298_ (
);

OR2X2 _11583_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_1607_)
);

DFFSR _11163_ (
    .CLK(clk_bF$buf54),
    .D(_1323_[30]),
    .Q(\datapath_1.regfile_1.regOut[21] [30]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL_0__17104_ (
);

DFFSR _9731_ (
    .CLK(clk_bF$buf109),
    .D(_597_[17]),
    .Q(\datapath_1.regfile_1.regOut[10] [17]),
    .R(rst_bF$buf84),
    .S(vdd)
);

FILL FILL65360x14820 (
);

AND2X2 _9311_ (
    .A(_452_),
    .B(_451_),
    .Y(_399_[26])
);

NOR2X1 _12788_ (
    .A(_2351_),
    .B(_2352_),
    .Y(_2353_)
);

AND2X2 _12368_ (
    .A(_2010_),
    .B(_2009_),
    .Y(_1983_[13])
);

FILL FILL_0__18729_ (
);

FILL FILL_0__18309_ (
);

FILL FILL_0__13864_ (
);

FILL FILL_0__13444_ (
);

FILL FILL446880x138320 (
);

FILL FILL491720x113620 (
);

FILL FILL400520x311220 (
);

FILL FILL_1__15236_ (
);

FILL FILL_1__10791_ (
);

OR2X2 _14934_ (
    .A(\datapath_1.mux_pcsrc.dout [16]),
    .B(_4001__bF$buf2),
    .Y(_3969_)
);

FILL FILL_0__14229_ (
);

OR2X2 _14514_ (
    .A(memoryOutData[5]),
    .B(_3803__bF$buf0),
    .Y(_3749_)
);

FILL FILL330600x316160 (
);

FILL FILL_0__18482_ (
);

FILL FILL232560x74100 (
);

FILL FILL_0__18062_ (
);

FILL FILL242440x281580 (
);

OR2X2 _15719_ (
    .A(_4669_),
    .B(_4666_),
    .Y(_4670_)
);

FILL FILL_0__10989_ (
);

OR2X2 _10854_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_1241_)
);

FILL FILL_0__10569_ (
);

OR2X2 _10434_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_1021_)
);

FILL FILL_0__10149_ (
);

OR2X2 _10014_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_801_)
);

FILL FILL448400x306280 (
);

FILL FILL_0__11510_ (
);

DFFSR _19552_ (
    .CLK(clk_bF$buf11),
    .D(_8320_[29]),
    .Q(\datapath_1.regfile_1.regOut[0] [29]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _19132_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_8031_)
);

FILL FILL434720x330980 (
);

FILL FILL_0__9788_ (
);

AND2X2 _11639_ (
    .A(_1644_),
    .B(_1643_),
    .Y(_1587_[28])
);

AND2X2 _11219_ (
    .A(_1424_),
    .B(_1423_),
    .Y(_1389_[17])
);

FILL FILL276640x24700 (
);

FILL FILL_1__13722_ (
);

FILL FILL_0__12715_ (
);

FILL FILL_1__16194_ (
);

AND2X2 _15892_ (
    .A(_4175__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_4840_)
);

FILL FILL253080x24700 (
);

AND2X2 _15472_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_4427_)
);

FILL FILL_0__15187_ (
);

AND2X2 _15052_ (
    .A(_4040_),
    .B(_4036_),
    .Y(_4041_)
);

FILL FILL77520x291460 (
);

FILL FILL464360x192660 (
);

FILL FILL182400x335920 (
);

AND2X2 _16677_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_5613_)
);

OR2X2 _16257_ (
    .A(_5198_),
    .B(_5195_),
    .Y(_5199_)
);

DFFSR _11392_ (
    .CLK(clk_bF$buf43),
    .D(_1455_[1]),
    .Q(\datapath_1.regfile_1.regOut[23] [1]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL_1__9109_ (
);

FILL FILL_0__17753_ (
);

FILL FILL_0__17333_ (
);

FILL FILL381520x296400 (
);

OR2X2 _8599_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .B(_134__bF$buf4),
    .Y(_78_)
);

FILL FILL_1__10427_ (
);

OR2X2 _9960_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_785_)
);

OR2X2 _9540_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_565_)
);

OR2X2 _9120_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [6]),
    .Y(_345_)
);

NAND2X1 _12597_ (
    .A(\datapath_1.alu_1.ALUInA [30]),
    .B(_2161_),
    .Y(_2162_)
);

DFFSR _12177_ (
    .CLK(clk_bF$buf103),
    .D(_1851_[12]),
    .Q(\datapath_1.regfile_1.regOut[29] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

FILL FILL_0__18958_ (
);

AND2X2 _18823_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_7727_)
);

FILL FILL_0__18538_ (
);

FILL FILL_0_BUFX2_insert400 (
);

FILL FILL_0_BUFX2_insert401 (
);

AND2X2 _18403_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_7313_)
);

FILL FILL_0_BUFX2_insert402 (
);

FILL FILL_0_BUFX2_insert403 (
);

FILL FILL_0_BUFX2_insert404 (
);

FILL FILL_0__13673_ (
);

FILL FILL_0_BUFX2_insert405 (
);

FILL FILL_0_BUFX2_insert407 (
);

FILL FILL_0_BUFX2_insert409 (
);

FILL FILL427120x326040 (
);

FILL FILL307800x276640 (
);

FILL FILL240160x330980 (
);

FILL FILL148960x217360 (
);

DFFSR _14743_ (
    .CLK(clk_bF$buf38),
    .D(_3804_[20]),
    .Q(\datapath_1.a [20]),
    .R(rst_bF$buf70),
    .S(vdd)
);

FILL FILL_0__14458_ (
);

FILL FILL_0__14038_ (
);

AND2X2 _14323_ (
    .A(_3661_),
    .B(_3660_),
    .Y(_3606_[27])
);

FILL FILL275120x237120 (
);

FILL FILL471200x93860 (
);

FILL FILL133000x74100 (
);

FILL FILL58520x103740 (
);

FILL FILL_0__18291_ (
);

OR2X2 _15948_ (
    .A(_4894_),
    .B(_4893_),
    .Y(_4895_)
);

OR2X2 _15528_ (
    .A(_4474_),
    .B(_4481_),
    .Y(_4482_)
);

AND2X2 _15108_ (
    .A(_4088_),
    .B(_4036_),
    .Y(_4089_)
);

FILL FILL_0__8392_ (
);

FILL FILL_0__10798_ (
);

OR2X2 _10663_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_1190__bF$buf2),
    .Y(_1134_)
);

FILL FILL_1__17611_ (
);

DFFSR _10243_ (
    .CLK(clk_bF$buf103),
    .D(_861_[13]),
    .Q(\datapath_1.regfile_1.regOut[14] [13]),
    .R(rst_bF$buf45),
    .S(vdd)
);

FILL FILL_0__16604_ (
);

AND2X2 _19361_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_8256_)
);

FILL FILL_0__19076_ (
);

FILL FILL75240x340860 (
);

DFFSR _8811_ (
    .CLK(clk_bF$buf96),
    .D(_135_[0]),
    .Q(\datapath_1.regfile_1.regOut[3] [0]),
    .R(rst_bF$buf72),
    .S(vdd)
);

FILL FILL493240x227240 (
);

FILL FILL_0__9177_ (
);

OR2X2 _11868_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_1757_)
);

OR2X2 _11448_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_1537_)
);

DFFSR _11028_ (
    .CLK(clk_bF$buf6),
    .D(_1257_[24]),
    .Q(\datapath_1.regfile_1.regOut[20] [24]),
    .R(rst_bF$buf31),
    .S(vdd)
);

FILL FILL_1__13111_ (
);

FILL FILL_0__17809_ (
);

FILL FILL_0__12944_ (
);

FILL FILL_0__12524_ (
);

AND2X2 _15281_ (
    .A(_4134_),
    .B(_4144_),
    .Y(_4239_)
);

FILL FILL419520x207480 (
);

FILL FILL_0__13729_ (
);

FILL FILL_0__13309_ (
);

FILL FILL191520x74100 (
);

OR2X2 _16486_ (
    .A(_5423_),
    .B(_5424_),
    .Y(_5425_)
);

FILL FILL136040x360620 (
);

AND2X2 _16066_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_5011_)
);

FILL FILL_0__17982_ (
);

FILL FILL_0__17562_ (
);

FILL FILL_0__17142_ (
);

FILL FILL322240x375440 (
);

FILL FILL113240x69160 (
);

FILL FILL468160x232180 (
);

FILL FILL_1__19354_ (
);

OR2X2 _18632_ (
    .A(_7537_),
    .B(_7538_),
    .Y(_7539_)
);

AND2X2 _18212_ (
    .A(_6317__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_7125_)
);

FILL FILL_0__13482_ (
);

FILL FILL_0__13062_ (
);

FILL FILL22800x345800 (
);

FILL FILL_0__8868_ (
);

OR2X2 _10719_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_1171_)
);

FILL FILL284240x355680 (
);

FILL FILL195320x74100 (
);

AND2X2 _19417_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_8312_)
);

FILL FILL_0__14687_ (
);

OR2X2 _14972_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.PCJump [29]),
    .Y(_3994_)
);

FILL FILL_0__14267_ (
);

OR2X2 _14552_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump [20]),
    .Y(_3774_)
);

AND2X2 _14132_ (
    .A(_3352__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3533_)
);

FILL FILL298680x316160 (
);

FILL FILL_1__16059_ (
);

AND2X2 _15757_ (
    .A(_4217__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_4707_)
);

FILL FILL233320x326040 (
);

AND2X2 _15337_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_4294_)
);

DFFSR _10892_ (
    .CLK(clk_bF$buf53),
    .D(_1191_[17]),
    .Q(\datapath_1.regfile_1.regOut[19] [17]),
    .R(rst_bF$buf111),
    .S(vdd)
);

AND2X2 _10472_ (
    .A(_1046_),
    .B(_1045_),
    .Y(_993_[26])
);

AND2X2 _10052_ (
    .A(_826_),
    .B(_825_),
    .Y(_795_[15])
);

FILL FILL_1__17000_ (
);

FILL FILL_0__16833_ (
);

FILL FILL12160x54340 (
);

FILL FILL392160x197600 (
);

AND2X2 _19170_ (
    .A(_6312__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .Y(_8068_)
);

FILL FILL415720x237120 (
);

OR2X2 _8620_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .B(_134__bF$buf4),
    .Y(_92_)
);

DFFSR _11677_ (
    .CLK(clk_bF$buf84),
    .D(_1587_[28]),
    .Q(\datapath_1.regfile_1.regOut[25] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL145920x251940 (
);

OR2X2 _11257_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_1454__bF$buf1),
    .Y(_1450_)
);

FILL FILL_1__13760_ (
);

FILL FILL_1__13340_ (
);

FILL FILL_0__17618_ (
);

OR2X2 _17903_ (
    .A(_6820_),
    .B(_6817_),
    .Y(_6821_)
);

FILL FILL_0__12333_ (
);

FILL FILL282720x311220 (
);

AND2X2 _15090_ (
    .A(_4074_),
    .B(_4073_),
    .Y(\datapath_1.regfile_1.regEn [5])
);

OR2X2 _9825_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_715_)
);

OR2X2 _9405_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_495_)
);

FILL FILL_1__8782_ (
);

FILL FILL269040x222300 (
);

FILL FILL193040x98800 (
);

FILL FILL201400x54340 (
);

FILL FILL_1__14545_ (
);

FILL FILL175560x69160 (
);

FILL FILL_0__13958_ (
);

OR2X2 _13823_ (
    .A(\datapath_1.a [2]),
    .B(_3342__bF$buf3),
    .Y(_3282_)
);

FILL FILL_0__13538_ (
);

INVX1 _13403_ (
    .A(_2930_),
    .Y(_2939_)
);

OR2X2 _16295_ (
    .A(_5233_),
    .B(_5236_),
    .Y(_5237_)
);

FILL FILL_0__17791_ (
);

FILL FILL63840x251940 (
);

FILL FILL_1__10045_ (
);

DFFSR _14608_ (
    .CLK(clk_bF$buf2),
    .D(_3738_[14]),
    .Q(\datapath_1.PCJump [16]),
    .R(rst_bF$buf33),
    .S(vdd)
);

FILL FILL297920x167960 (
);

FILL FILL_0__18576_ (
);

AND2X2 _18861_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_7764_)
);

FILL FILL_0__18156_ (
);

OR2X2 _18441_ (
    .A(_7349_),
    .B(_7350_),
    .Y(_7351_)
);

OR2X2 _18021_ (
    .A(_6936_),
    .B(_6935_),
    .Y(_6937_)
);

FILL FILL_0__13291_ (
);

FILL FILL179360x69160 (
);

FILL FILL_0__8677_ (
);

OR2X2 _10948_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_1322__bF$buf0),
    .Y(_1284_)
);

OR2X2 _10528_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_1124__bF$buf4),
    .Y(_1064_)
);

DFFSR _10108_ (
    .CLK(clk_bF$buf39),
    .D(_795_[7]),
    .Q(\datapath_1.regfile_1.regOut[13] [7]),
    .R(rst_bF$buf80),
    .S(vdd)
);

OR2X2 _19226_ (
    .A(_8123_),
    .B(_8116_),
    .Y(_8124_)
);

OR2X2 _14781_ (
    .A(\datapath_1.rd2 [8]),
    .B(_3935__bF$buf3),
    .Y(_3887_)
);

DFFSR _14361_ (
    .CLK(clk_bF$buf12),
    .D(_3606_[25]),
    .Q(ALUOut[25]),
    .R(rst_bF$buf91),
    .S(vdd)
);

FILL FILL174040x326040 (
);

FILL FILL291840x242060 (
);

FILL FILL_0__12809_ (
);

FILL FILL160360x350740 (
);

FILL FILL_1__16288_ (
);

OR2X2 _15986_ (
    .A(_4931_),
    .B(_4932_),
    .Y(_4933_)
);

AND2X2 _15566_ (
    .A(_4135__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_4519_)
);

AOI22X1 _15146_ (
    .A(\datapath_1.a3 [4]),
    .B(_4024_),
    .C(_4020_),
    .D(_4054_),
    .Y(_4113_)
);

FILL FILL227240x64220 (
);

OR2X2 _10281_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_939_)
);

FILL FILL8360x158080 (
);

FILL FILL278920x113620 (
);

FILL FILL_0__16222_ (
);

FILL FILL164160x271700 (
);

AND2X2 _11486_ (
    .A(_1562_),
    .B(_1561_),
    .Y(_1521_[20])
);

AND2X2 _11066_ (
    .A(_1342_),
    .B(_1341_),
    .Y(_1323_[9])
);

FILL FILL101080x202540 (
);

FILL FILL_0__17847_ (
);

FILL FILL117800x316160 (
);

FILL FILL_0__17427_ (
);

AND2X2 _17712_ (
    .A(_6236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_6633_)
);

FILL FILL_0__17007_ (
);

FILL FILL_0__12982_ (
);

FILL FILL_0__12562_ (
);

FILL FILL_0__12142_ (
);

FILL FILL190760x39520 (
);

OR2X2 _9634_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .B(_662__bF$buf1),
    .Y(_608_)
);

DFFSR _9214_ (
    .CLK(clk_bF$buf107),
    .D(_333_[16]),
    .Q(\datapath_1.regfile_1.regOut[6] [16]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL_1__8591_ (
);

FILL FILL382280x261820 (
);

FILL FILL_1__19219_ (
);

FILL FILL381520x0 (
);

AND2X2 _18917_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_7819_)
);

FILL FILL_0__13767_ (
);

FILL FILL_0__13347_ (
);

OR2X2 _13632_ (
    .A(_3121_),
    .B(_3118_),
    .Y(\datapath_1.mux_pcsrc.dout [5])
);

XOR2X1 _13212_ (
    .A(_2212_),
    .B(_2746_),
    .Y(_2760_)
);

FILL FILL_1__9796_ (
);

FILL FILL_0__17180_ (
);

OR2X2 _14837_ (
    .A(vdd),
    .B(_2_[27]),
    .Y(_3924_)
);

OR2X2 _14417_ (
    .A(vdd),
    .B(\datapath_1.Data [16]),
    .Y(_3704_)
);

FILL FILL_1__16500_ (
);

FILL FILL339720x227240 (
);

AND2X2 _18670_ (
    .A(_6229__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_7576_)
);

OR2X2 _18250_ (
    .A(_7159_),
    .B(_7162_),
    .Y(_7163_)
);

FILL FILL_1__11479_ (
);

FILL FILL225720x345800 (
);

FILL FILL114000x163020 (
);

DFFSR _10757_ (
    .CLK(clk_bF$buf73),
    .D(_1125_[11]),
    .Q(\datapath_1.regfile_1.regOut[18] [11]),
    .R(rst_bF$buf39),
    .S(vdd)
);

AND2X2 _10337_ (
    .A(_976_),
    .B(_975_),
    .Y(_927_[24])
);

FILL FILL_1__12840_ (
);

FILL FILL443840x148200 (
);

FILL FILL_0__11833_ (
);

OR2X2 _19455_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8339_)
);

AND2X2 _19035_ (
    .A(_7935_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd1 [25])
);

AND2X2 _14590_ (
    .A(_3799_),
    .B(_3798_),
    .Y(_3738_[30])
);

OR2X2 _14170_ (
    .A(MemToReg_bF$buf1),
    .B(ALUOut[9]),
    .Y(_3558_)
);

OR2X2 _8905_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .B(_266__bF$buf4),
    .Y(_242_)
);

FILL FILL289560x64220 (
);

FILL FILL473480x64220 (
);

FILL FILL84360x207480 (
);

FILL FILL_1__13205_ (
);

AOI21X1 _12903_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .B(\datapath_1.alu_1.ALUInB [20]),
    .C(_2467_),
    .Y(_2468_)
);

FILL FILL_1_BUFX2_insert333 (
);

FILL FILL_1_BUFX2_insert335 (
);

FILL FILL_1_BUFX2_insert337 (
);

AND2X2 _15795_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_4745_)
);

OR2X2 _15375_ (
    .A(_4329_),
    .B(_4330_),
    .Y(_4331_)
);

OR2X2 _10090_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .B(_860__bF$buf0),
    .Y(_852_)
);

FILL FILL_0__16871_ (
);

FILL FILL_0__16451_ (
);

FILL FILL_0__16031_ (
);

FILL FILL51680x9880 (
);

FILL FILL300960x350740 (
);

INVX2 _11295_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .Y(_1520_)
);

FILL FILL38760x19760 (
);

AND2X2 _17941_ (
    .A(_6312__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_6858_)
);

FILL FILL_0__17656_ (
);

OR2X2 _17521_ (
    .A(_6437_),
    .B(_6444_),
    .Y(_6445_)
);

AND2X2 _17101_ (
    .A(_4228__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_6030_)
);

FILL FILL_0__12791_ (
);

FILL FILL_0__12371_ (
);

DFFSR _9863_ (
    .CLK(clk_bF$buf46),
    .D(_663_[20]),
    .Q(\datapath_1.regfile_1.regOut[11] [20]),
    .R(rst_bF$buf57),
    .S(vdd)
);

AND2X2 _9443_ (
    .A(_520_),
    .B(_519_),
    .Y(_465_[27])
);

AND2X2 _9023_ (
    .A(_300_),
    .B(_299_),
    .Y(_267_[16])
);

FILL FILL152000x197600 (
);

FILL FILL_1__19448_ (
);

FILL FILL_1__14163_ (
);

OR2X2 _18726_ (
    .A(_7623_),
    .B(_7630_),
    .Y(_7631_)
);

AND2X2 _18306_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_7218_)
);

FILL FILL_0__13996_ (
);

FILL FILL383800x182780 (
);

OR2X2 _13861_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [15]),
    .Y(_3307_)
);

FILL FILL_0__13156_ (
);

AND2X2 _13441_ (
    .A(_2623_),
    .B(_2528_),
    .Y(_2974_)
);

NOR3X1 _13021_ (
    .A(_2579_),
    .B(_2576_),
    .C(_2577_),
    .Y(_2580_)
);

FILL FILL5320x192660 (
);

FILL FILL_0__9903_ (
);

FILL FILL_1__15788_ (
);

FILL FILL315400x143260 (
);

OR2X2 _14646_ (
    .A(\datapath_1.rd1 [6]),
    .B(_3869__bF$buf0),
    .Y(_3817_)
);

AND2X2 _14226_ (
    .A(_3595_),
    .B(_3594_),
    .Y(\datapath_1.mux_wd3.dout [27])
);

FILL FILL_0__15722_ (
);

FILL FILL_0__15302_ (
);

FILL FILL_0__18194_ (
);

FILL FILL251560x0 (
);

OR2X2 _10986_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_1309_)
);

OR2X2 _10566_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_1089_)
);

OR2X2 _10146_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_869_)
);

FILL FILL_0__16927_ (
);

FILL FILL_0__11642_ (
);

FILL FILL_0__11222_ (
);

FILL FILL_0__19399_ (
);

OR2X2 _19264_ (
    .A(_8159_),
    .B(_8160_),
    .Y(_8161_)
);

OR2X2 _8714_ (
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .Y(_199_)
);

FILL FILL241680x163020 (
);

FILL FILL_1__13854_ (
);

FILL FILL505400x266760 (
);

FILL FILL_0__12847_ (
);

XNOR2X1 _12712_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2277_)
);

AND2X2 _15184_ (
    .A(_4141_),
    .B(_4139_),
    .Y(_4142_)
);

OR2X2 _9919_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .B(_794__bF$buf2),
    .Y(_758_)
);

FILL FILL433960x212420 (
);

FILL FILL213560x296400 (
);

FILL FILL_0__16680_ (
);

FILL FILL262960x19760 (
);

FILL FILL_0__16260_ (
);

FILL FILL281200x138320 (
);

AND2X2 _13917_ (
    .A(_3347__bF$buf2),
    .B(\aluControl_1.inst [0]),
    .Y(_3348_)
);

FILL FILL350360x59280 (
);

FILL FILL177080x108680 (
);

AND2X2 _16389_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_5329_)
);

FILL FILL376960x163020 (
);

FILL FILL_1__18472_ (
);

FILL FILL_1__18052_ (
);

OR2X2 _17750_ (
    .A(_6665_),
    .B(_6669_),
    .Y(_6670_)
);

FILL FILL_0__17045_ (
);

AND2X2 _17330_ (
    .A(_6255__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_6256_)
);

FILL FILL_1__10139_ (
);

OR2X2 _9672_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_633_)
);

OR2X2 _9252_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_413_)
);

FILL FILL_1__11500_ (
);

FILL FILL_0__10913_ (
);

FILL FILL377720x59280 (
);

INVX1 _18955_ (
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_7857_)
);

OR2X2 _18535_ (
    .A(_7441_),
    .B(_7442_),
    .Y(_7443_)
);

AND2X2 _18115_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_7030_)
);

FILL FILL_0__13385_ (
);

OR2X2 _13670_ (
    .A(_3152_),
    .B(_3153_),
    .Y(_3154_)
);

OR2X2 _13250_ (
    .A(_2157__bF$buf3),
    .B(_2794_),
    .Y(_2795_)
);

FILL FILL110200x286520 (
);

FILL FILL399760x113620 (
);

FILL FILL424840x83980 (
);

FILL FILL103360x14820 (
);

FILL FILL107160x237120 (
);

FILL FILL_1__12705_ (
);

FILL FILL106400x79040 (
);

FILL FILL123120x29640 (
);

FILL FILL_1__15177_ (
);

DFFSR _14875_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[23]),
    .Q(_2_[23]),
    .R(rst_bF$buf61),
    .S(vdd)
);

AND2X2 _14455_ (
    .A(_3729_),
    .B(_3728_),
    .Y(_3672_[28])
);

OR2X2 _14035_ (
    .A(_3449_),
    .B(_3448_),
    .Y(_3450_)
);

FILL FILL41800x281580 (
);

FILL FILL238640x316160 (
);

FILL FILL_0__15951_ (
);

FILL FILL228000x276640 (
);

FILL FILL345800x192660 (
);

FILL FILL224960x340860 (
);

OR2X2 _10795_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .B(_1256__bF$buf0),
    .Y(_1202_)
);

DFFSR _10375_ (
    .CLK(clk_bF$buf5),
    .D(_927_[16]),
    .Q(\datapath_1.regfile_1.regOut[15] [16]),
    .R(rst_bF$buf10),
    .S(vdd)
);

FILL FILL_0__16736_ (
);

OR2X2 _16601_ (
    .A(_5522_),
    .B(_5537_),
    .Y(_5538_)
);

FILL FILL_0__16316_ (
);

FILL FILL_0__11871_ (
);

FILL FILL_0__11451_ (
);

FILL FILL332120x197600 (
);

OR2X2 _19493_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_8364_)
);

OR2X2 _19073_ (
    .A(_7969_),
    .B(_7972_),
    .Y(_7973_)
);

FILL FILL259920x247000 (
);

FILL FILL281200x365560 (
);

DFFSR _8943_ (
    .CLK(clk_bF$buf44),
    .D(_201_[3]),
    .Q(\datapath_1.regfile_1.regOut[4] [3]),
    .R(rst_bF$buf97),
    .S(vdd)
);

OR2X2 _8523_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_47_)
);

FILL FILL365560x321100 (
);

FILL FILL_1__18948_ (
);

FILL FILL254600x44460 (
);

AND2X2 _17806_ (
    .A(_6328__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_6725_)
);

NAND2X1 _12941_ (
    .A(_2504_),
    .B(_2167_),
    .Y(_2505_)
);

FILL FILL_0__12656_ (
);

FILL FILL_1_BUFX2_insert713 (
);

OR2X2 _12521_ (
    .A(\control_1.op [4]),
    .B(\control_1.op [5]),
    .Y(_2111_)
);

AND2X2 _12101_ (
    .A(_1872_),
    .B(_1871_),
    .Y(_1851_[10])
);

FILL FILL_1_BUFX2_insert715 (
);

FILL FILL_1_BUFX2_insert717 (
);

FILL FILL231040x44460 (
);

DFFSR _9728_ (
    .CLK(clk_bF$buf13),
    .D(_597_[14]),
    .Q(\datapath_1.regfile_1.regOut[10] [14]),
    .R(rst_bF$buf90),
    .S(vdd)
);

AND2X2 _9308_ (
    .A(_450_),
    .B(_449_),
    .Y(_399_[25])
);

FILL FILL303240x281580 (
);

FILL FILL294120x177840 (
);

FILL FILL102600x167960 (
);

FILL FILL_1__14028_ (
);

FILL FILL376960x256880 (
);

OR2X2 _13726_ (
    .A(_3200_),
    .B(_3201_),
    .Y(_3202_)
);

INVX1 _13306_ (
    .A(_2847_),
    .Y(\datapath_1.ALUResult [8])
);

FILL FILL114000x83980 (
);

AND2X2 _16198_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_5141_)
);

FILL FILL_0__17694_ (
);

FILL FILL_0__17274_ (
);

FILL FILL53200x306280 (
);

DFFSR _9481_ (
    .CLK(clk_bF$buf60),
    .D(_465_[25]),
    .Q(\datapath_1.regfile_1.regOut[8] [25]),
    .R(rst_bF$buf101),
    .S(vdd)
);

OR2X2 _9061_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .B(_332__bF$buf2),
    .Y(_326_)
);

FILL FILL357200x217360 (
);

FILL FILL_0__10722_ (
);

FILL FILL_0__10302_ (
);

FILL FILL_0__18899_ (
);

AND2X2 _18764_ (
    .A(_6293__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_7669_)
);

FILL FILL386080x345800 (
);

OR2X2 _18344_ (
    .A(_7254_),
    .B(_7253_),
    .Y(_7255_)
);

FILL FILL_0__18059_ (
);

FILL FILL_0__19420_ (
);

FILL FILL429400x256880 (
);

FILL FILL275120x123500 (
);

FILL FILL_0__9521_ (
);

FILL FILL_0__9101_ (
);

FILL FILL_0__11507_ (
);

FILL FILL461320x138320 (
);

DFFSR _19549_ (
    .CLK(clk_bF$buf86),
    .D(_8320_[26]),
    .Q(\datapath_1.regfile_1.regOut[0] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

OR2X2 _19129_ (
    .A(_8027_),
    .B(_8014_),
    .Y(_8028_)
);

OR2X2 _14684_ (
    .A(vdd),
    .B(\datapath_1.a [19]),
    .Y(_3842_)
);

FILL FILL_0__14399_ (
);

OR2X2 _14264_ (
    .A(vdd),
    .B(ALUOut[8]),
    .Y(_3622_)
);

FILL FILL15960x286520 (
);

FILL FILL60800x261820 (
);

FILL FILL464360x54340 (
);

FILL FILL_0__15340_ (
);

FILL FILL439280x247000 (
);

FILL FILL40280x64220 (
);

FILL FILL100320x350740 (
);

FILL FILL51680x365560 (
);

AND2X2 _15889_ (
    .A(_4154__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_4837_)
);

AND2X2 _15469_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_4424_)
);

AND2X2 _15049_ (
    .A(_4031_),
    .B(_4018_),
    .Y(_4038_)
);

AND2X2 _10184_ (
    .A(_894_),
    .B(_893_),
    .Y(_861_[16])
);

FILL FILL_0__16965_ (
);

FILL FILL_0__16545_ (
);

AND2X2 _16830_ (
    .A(_4197__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_5763_)
);

AND2X2 _16410_ (
    .A(_4175__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_5350_)
);

FILL FILL_0__16125_ (
);

FILL FILL_0__11260_ (
);

OR2X2 _8752_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .B(_200__bF$buf4),
    .Y(_160_)
);

FILL FILL12920x182780 (
);

OR2X2 _11389_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .B(_1520__bF$buf4),
    .Y(_1518_)
);

FILL FILL_1__18337_ (
);

OR2X2 _17615_ (
    .A(_6535_),
    .B(_6536_),
    .Y(_6537_)
);

FILL FILL_0__12885_ (
);

AND2X2 _12750_ (
    .A(_2309_),
    .B(_2314_),
    .Y(_2315_)
);

OR2X2 _12330_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_1985_)
);

OR2X2 _9957_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_783_)
);

OR2X2 _9537_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_563_)
);

OR2X2 _9117_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_343_)
);

FILL FILL421040x24700 (
);

FILL FILL_1__8494_ (
);

FILL FILL_1__14677_ (
);

FILL FILL_0_BUFX2_insert370 (
);

FILL FILL_0_BUFX2_insert372 (
);

FILL FILL_0_BUFX2_insert374 (
);

OR2X2 _13955_ (
    .A(_3379_),
    .B(_3380_),
    .Y(_3381_)
);

OR2X2 _13535_ (
    .A(ALUOut[15]),
    .B(_3079__bF$buf0),
    .Y(_3045_)
);

OR2X2 _13115_ (
    .A(_2288_),
    .B(_2667_),
    .Y(_2668_)
);

FILL FILL_0_BUFX2_insert376 (
);

FILL FILL_0_BUFX2_insert377 (
);

FILL FILL_0_BUFX2_insert378 (
);

FILL FILL_0_BUFX2_insert379 (
);

FILL FILL22040x271700 (
);

FILL FILL61560x88920 (
);

FILL FILL_1__18090_ (
);

FILL FILL_1__10177_ (
);

AND2X2 _9290_ (
    .A(_438_),
    .B(_437_),
    .Y(_399_[19])
);

FILL FILL135280x335920 (
);

FILL FILL_0__15816_ (
);

FILL FILL_0__10951_ (
);

FILL FILL_0__10531_ (
);

OR2X2 _18993_ (
    .A(_7893_),
    .B(_7892_),
    .Y(_7894_)
);

FILL FILL_0__18288_ (
);

AND2X2 _18573_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_7481_)
);

OR2X2 _18153_ (
    .A(_7066_),
    .B(_7059_),
    .Y(_7067_)
);

FILL FILL152760x345800 (
);

FILL FILL402800x311220 (
);

FILL FILL_0__11316_ (
);

OR2X2 _11601_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_1619_)
);

FILL FILL462840x74100 (
);

OR2X2 _19358_ (
    .A(_8222_),
    .B(_8253_),
    .Y(_8254_)
);

FILL FILL233320x212420 (
);

DFFSR _14493_ (
    .CLK(clk_bF$buf42),
    .D(_3672_[28]),
    .Q(\datapath_1.Data [28]),
    .R(rst_bF$buf100),
    .S(vdd)
);

AND2X2 _14073_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3482_)
);

OR2X2 _8808_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_197_)
);

FILL FILL500840x291460 (
);

FILL FILL244720x281580 (
);

FILL FILL205960x247000 (
);

FILL FILL_1__13528_ (
);

AND2X2 _12806_ (
    .A(_2370_),
    .B(_2162_),
    .Y(_2371_)
);

AND2X2 _15698_ (
    .A(_4197__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_4649_)
);

AND2X2 _15278_ (
    .A(_4129_),
    .B(_4144_),
    .Y(_4236_)
);

FILL FILL28120x128440 (
);

FILL FILL_0__16774_ (
);

FILL FILL_1__9911_ (
);

AND2X2 _8981_ (
    .A(_272_),
    .B(_271_),
    .Y(_267_[2])
);

DFFSR _8561_ (
    .CLK(clk_bF$buf91),
    .D(_3_[8]),
    .Q(\datapath_1.regfile_1.regOut[1] [8]),
    .R(rst_bF$buf74),
    .S(vdd)
);

FILL FILL_1__18986_ (
);

FILL FILL_1__18566_ (
);

AND2X2 _11198_ (
    .A(_1410_),
    .B(_1409_),
    .Y(_1389_[10])
);

FILL FILL245480x247000 (
);

FILL FILL_1__13281_ (
);

FILL FILL_0__17559_ (
);

OR2X2 _17844_ (
    .A(_6761_),
    .B(_6762_),
    .Y(_6763_)
);

FILL FILL455240x123500 (
);

OR2X2 _17424_ (
    .A(_6348_),
    .B(_6345_),
    .Y(_6349_)
);

FILL FILL_0__17139_ (
);

AND2X2 _17004_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_5935_)
);

FILL FILL_0__12274_ (
);

FILL FILL_0__18500_ (
);

FILL FILL94240x163020 (
);

OR2X2 _9766_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_728__bF$buf2),
    .Y(_676_)
);

DFFSR _9346_ (
    .CLK(clk_bF$buf81),
    .D(_399_[19]),
    .Q(\datapath_1.regfile_1.regOut[7] [19]),
    .R(rst_bF$buf101),
    .S(vdd)
);

FILL FILL440800x345800 (
);

FILL FILL_0__8601_ (
);

OR2X2 _18629_ (
    .A(_7535_),
    .B(_7534_),
    .Y(_7536_)
);

OR2X2 _18209_ (
    .A(_7120_),
    .B(_7121_),
    .Y(_7122_)
);

FILL FILL_0__13899_ (
);

FILL FILL_0__13479_ (
);

OR2X2 _13764_ (
    .A(_3234_),
    .B(_3233_),
    .Y(_3235_)
);

FILL FILL325280x34580 (
);

MUX2X1 _13344_ (
    .A(_2376__bF$buf1),
    .B(_2883_),
    .S(_2882_),
    .Y(_2884_)
);

FILL FILL_0__14840_ (
);

FILL FILL_0__14420_ (
);

FILL FILL_0__9806_ (
);

OR2X2 _14969_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.PCJump [28]),
    .Y(_3992_)
);

OR2X2 _14549_ (
    .A(IRWrite_bF$buf0),
    .B(\datapath_1.PCJump [19]),
    .Y(_3772_)
);

AND2X2 _14129_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3530_)
);

OR2X2 _15910_ (
    .A(_4857_),
    .B(_4856_),
    .Y(_4858_)
);

FILL FILL_0__15205_ (
);

FILL FILL_0__10340_ (
);

FILL FILL_0__18097_ (
);

OR2X2 _18382_ (
    .A(_7292_),
    .B(_7277_),
    .Y(_7293_)
);

FILL FILL415720x350740 (
);

DFFSR _10889_ (
    .CLK(clk_bF$buf98),
    .D(_1191_[14]),
    .Q(\datapath_1.regfile_1.regOut[19] [14]),
    .R(rst_bF$buf87),
    .S(vdd)
);

FILL FILL_1__17417_ (
);

AND2X2 _10469_ (
    .A(_1044_),
    .B(_1043_),
    .Y(_993_[25])
);

AND2X2 _10049_ (
    .A(_824_),
    .B(_823_),
    .Y(_795_[14])
);

FILL FILL_1__12972_ (
);

FILL FILL_1__12552_ (
);

FILL FILL_0__11965_ (
);

OR2X2 _11830_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .B(_1784__bF$buf1),
    .Y(_1732_)
);

FILL FILL345800x355680 (
);

DFFSR _11410_ (
    .CLK(clk_bF$buf19),
    .D(_1455_[19]),
    .Q(\datapath_1.regfile_1.regOut[23] [19]),
    .R(rst_bF$buf19),
    .S(vdd)
);

AND2X2 _19167_ (
    .A(_6216__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_8065_)
);

OR2X2 _8617_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .B(_134__bF$buf3),
    .Y(_90_)
);

OR2X2 _12615_ (
    .A(_2177_),
    .B(_2179_),
    .Y(_2180_)
);

AND2X2 _15087_ (
    .A(_4071_),
    .B(_4066_),
    .Y(_4072_)
);

FILL FILL_1__17590_ (
);

FILL FILL_1__17170_ (
);

FILL FILL112480x54340 (
);

FILL FILL_0__16163_ (
);

FILL FILL77520x340860 (
);

FILL FILL_1__9300_ (
);

FILL FILL117040x108680 (
);

OR2X2 _8790_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_185_)
);

FILL FILL12160x158080 (
);

FILL FILL_0__17788_ (
);

AND2X2 _17653_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_6575_)
);

FILL FILL_0__17368_ (
);

AND2X2 _17233_ (
    .A(_4167__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_6160_)
);

FILL FILL307040x79040 (
);

FILL FILL_0__12083_ (
);

DFFSR _9995_ (
    .CLK(clk_bF$buf101),
    .D(_729_[23]),
    .Q(\datapath_1.regfile_1.regOut[12] [23]),
    .R(rst_bF$buf54),
    .S(vdd)
);

AND2X2 _9575_ (
    .A(_588_),
    .B(_587_),
    .Y(_531_[28])
);

AND2X2 _9155_ (
    .A(_368_),
    .B(_367_),
    .Y(_333_[17])
);

FILL FILL_0__8410_ (
);

FILL FILL_1__14295_ (
);

AND2X2 _18858_ (
    .A(_6262__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_7761_)
);

FILL FILL_0_BUFX2_insert750 (
);

OR2X2 _18438_ (
    .A(_7347_),
    .B(_7344_),
    .Y(_7348_)
);

FILL FILL_0_BUFX2_insert752 (
);

OR2X2 _18018_ (
    .A(_6933_),
    .B(_6932_),
    .Y(_6934_)
);

OR2X2 _13993_ (
    .A(_3413_),
    .B(_3412_),
    .Y(_3414_)
);

FILL FILL_0_BUFX2_insert754 (
);

FILL FILL183160x143260 (
);

FILL FILL_0__13288_ (
);

OR2X2 _13573_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.PCJump [28]),
    .Y(_3070_)
);

INVX1 _13153_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .Y(_2704_)
);

FILL FILL_0_BUFX2_insert756 (
);

FILL FILL_0_BUFX2_insert757 (
);

FILL FILL_0_BUFX2_insert758 (
);

FILL FILL_0_BUFX2_insert759 (
);

FILL FILL324520x375440 (
);

OR2X2 _14778_ (
    .A(\datapath_1.rd2 [7]),
    .B(_3935__bF$buf0),
    .Y(_3885_)
);

DFFSR _14358_ (
    .CLK(clk_bF$buf12),
    .D(_3606_[22]),
    .Q(ALUOut[22]),
    .R(rst_bF$buf91),
    .S(vdd)
);

FILL FILL_0__15854_ (
);

FILL FILL_0__15434_ (
);

FILL FILL_0__15014_ (
);

FILL FILL172520x286520 (
);

AND2X2 _18191_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_7104_)
);

FILL FILL126920x133380 (
);

FILL FILL443080x261820 (
);

OR2X2 _10698_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_1157_)
);

FILL FILL459800x375440 (
);

OR2X2 _10278_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_937_)
);

FILL FILL_1__12361_ (
);

FILL FILL_0__16639_ (
);

OR2X2 _16924_ (
    .A(_5855_),
    .B(_5854_),
    .Y(_5856_)
);

OR2X2 _16504_ (
    .A(_5442_),
    .B(_5427_),
    .Y(_5443_)
);

FILL FILL_0__11774_ (
);

FILL FILL_0__11354_ (
);

AND2X2 _19396_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_8291_)
);

AND2X2 _8846_ (
    .A(_202_),
    .B(_265_),
    .Y(_201_[0])
);

FILL FILL218120x316160 (
);

BUFX2 _8426_ (
    .A(_2_[2]),
    .Y(memoryWriteData[2])
);

FILL FILL_1__13146_ (
);

AND2X2 _17709_ (
    .A(_6302__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_6630_)
);

FILL FILL_0__12979_ (
);

OR2X2 _12844_ (
    .A(_2401_),
    .B(_2408_),
    .Y(_2409_)
);

FILL FILL_0__12559_ (
);

FILL FILL220400x54340 (
);

DFFSR _12424_ (
    .CLK(clk_bF$buf4),
    .D(_1983_[1]),
    .Q(\datapath_1.regfile_1.regOut[31] [1]),
    .R(rst_bF$buf71),
    .S(vdd)
);

OR2X2 _12004_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .B(_1850__bF$buf1),
    .Y(_1828_)
);

FILL FILL136040x222300 (
);

FILL FILL_0__13920_ (
);

FILL FILL11400x24700 (
);

FILL FILL_0__16392_ (
);

AND2X2 _13629_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [5]),
    .Y(_3119_)
);

OAI21X1 _13209_ (
    .A(_2212_),
    .B(_2503_),
    .C(_2756_),
    .Y(_2757_)
);

FILL FILL_1__15712_ (
);

FILL FILL504640x148200 (
);

FILL FILL_0__14705_ (
);

FILL FILL403560x167960 (
);

AND2X2 _17882_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_6800_)
);

OR2X2 _17462_ (
    .A(_6386_),
    .B(_6385_),
    .Y(_6387_)
);

FILL FILL_0__17177_ (
);

AND2X2 _17042_ (
    .A(_4241__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_5972_)
);

FILL FILL284240x217360 (
);

OR2X2 _9384_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_481_)
);

FILL FILL_1__11632_ (
);

FILL FILL_1__19389_ (
);

AND2X2 _10910_ (
    .A(_1258_),
    .B(_1321_),
    .Y(_1257_[0])
);

AND2X2 _18667_ (
    .A(_6236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_7573_)
);

AND2X2 _18247_ (
    .A(_6323__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_7160_)
);

FILL FILL_0__13097_ (
);

OR2X2 _13382_ (
    .A(_2182_),
    .B(_2181_),
    .Y(_2919_)
);

FILL FILL_0__19323_ (
);

FILL FILL269040x296400 (
);

FILL FILL_0__9424_ (
);

AND2X2 _14587_ (
    .A(_3797_),
    .B(_3796_),
    .Y(_3738_[29])
);

OR2X2 _14167_ (
    .A(MemToReg_bF$buf1),
    .B(ALUOut[8]),
    .Y(_3556_)
);

FILL FILL4560x167960 (
);

FILL FILL_1__16670_ (
);

FILL FILL_0__15663_ (
);

FILL FILL_0__15243_ (
);

FILL FILL122360x256880 (
);

FILL FILL_1__17455_ (
);

FILL FILL_1__17035_ (
);

OR2X2 _10087_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .B(_860__bF$buf3),
    .Y(_850_)
);

AND2X2 _16733_ (
    .A(_4195__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_5668_)
);

FILL FILL_0__16028_ (
);

OR2X2 _16313_ (
    .A(_5254_),
    .B(_5223_),
    .Y(_5255_)
);

FILL FILL126920x271700 (
);

FILL FILL_0__11583_ (
);

FILL FILL176320x326040 (
);

OR2X2 _8655_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_115_)
);

FILL FILL162640x350740 (
);

FILL FILL_1__13795_ (
);

AND2X2 _17938_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_6855_)
);

AND2X2 _17518_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_6442_)
);

FILL FILL50160x24700 (
);

FILL FILL_0__12368_ (
);

XNOR2X1 _12653_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2218_)
);

AND2X2 _12233_ (
    .A(_1940_),
    .B(_1939_),
    .Y(_1917_[11])
);

FILL FILL142120x93860 (
);

FILL FILL_0_BUFX2_insert1100 (
);

FILL FILL63840x113620 (
);

FILL FILL_0_BUFX2_insert1101 (
);

FILL FILL40280x256880 (
);

FILL FILL_0_BUFX2_insert1102 (
);

FILL FILL_0_BUFX2_insert1103 (
);

FILL FILL490200x123500 (
);

FILL FILL_0_BUFX2_insert1105 (
);

FILL FILL_0_BUFX2_insert1107 (
);

FILL FILL_0_BUFX2_insert1109 (
);

OR2X2 _13858_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [14]),
    .Y(_3305_)
);

AND2X2 _13438_ (
    .A(_2971_),
    .B(_2968_),
    .Y(_2972_)
);

NOR2X1 _13018_ (
    .A(_2327_),
    .B(_2498_),
    .Y(_2577_)
);

FILL FILL103360x202540 (
);

FILL FILL286520x54340 (
);

FILL FILL380760x340860 (
);

FILL FILL_0__14514_ (
);

FILL FILL361760x177840 (
);

OR2X2 _17691_ (
    .A(_6608_),
    .B(_6611_),
    .Y(_6612_)
);

OR2X2 _17271_ (
    .A(_6190_),
    .B(_6197_),
    .Y(_6198_)
);

FILL FILL490200x69160 (
);

FILL FILL398240x237120 (
);

OR2X2 _9193_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .B(_398__bF$buf3),
    .Y(_394_)
);

FILL FILL_1__11441_ (
);

FILL FILL_0__15719_ (
);

FILL FILL_0__10854_ (
);

OR2X2 _18896_ (
    .A(_7797_),
    .B(_7798_),
    .Y(_7799_)
);

AND2X2 _18476_ (
    .A(_6250__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_7385_)
);

OR2X2 _18056_ (
    .A(_6964_),
    .B(_6971_),
    .Y(_6972_)
);

NAND2X1 _13191_ (
    .A(_2501_),
    .B(_2739_),
    .Y(_2740_)
);

FILL FILL433200x340860 (
);

FILL FILL_1__12646_ (
);

FILL FILL_0__9653_ (
);

FILL FILL_0__11639_ (
);

FILL FILL_0__9233_ (
);

DFFSR _11924_ (
    .CLK(clk_bF$buf6),
    .D(_1719_[17]),
    .Q(\datapath_1.regfile_1.regOut[27] [17]),
    .R(rst_bF$buf31),
    .S(vdd)
);

AND2X2 _11504_ (
    .A(_1574_),
    .B(_1573_),
    .Y(_1521_[26])
);

FILL FILL_0__11219_ (
);

OR2X2 _14396_ (
    .A(vdd),
    .B(\datapath_1.Data [9]),
    .Y(_3690_)
);

FILL FILL141360x370500 (
);

FILL FILL376200x291460 (
);

FILL FILL_0__15892_ (
);

AND2X2 _12709_ (
    .A(_2273_),
    .B(_2270_),
    .Y(_2274_)
);

FILL FILL_1__17684_ (
);

FILL FILL259160x360620 (
);

FILL FILL_0__16677_ (
);

AND2X2 _16962_ (
    .A(_4189__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_5893_)
);

AND2X2 _16542_ (
    .A(_4241__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_5480_)
);

FILL FILL_0__16257_ (
);

AND2X2 _16122_ (
    .A(_5066_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd2 [13])
);

FILL FILL86640x207480 (
);

FILL FILL189240x365560 (
);

OR2X2 _8884_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .B(_266__bF$buf2),
    .Y(_228_)
);

OR2X2 _8464_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .B(_68__bF$buf2),
    .Y(_8_)
);

FILL FILL_1__10712_ (
);

FILL FILL350360x335920 (
);

NOR2X1 _17747_ (
    .A(_6310__bF$buf4),
    .B(_6666_),
    .Y(_6667_)
);

OR2X2 _17327_ (
    .A(_6245_),
    .B(_6252_),
    .Y(_6253_)
);

FILL FILL_0__12597_ (
);

AND2X2 _12882_ (
    .A(_2444_),
    .B(_2446_),
    .Y(_2447_)
);

OR2X2 _12462_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2056_)
);

DFFSR _12042_ (
    .CLK(clk_bF$buf36),
    .D(_1785_[6]),
    .Q(\datapath_1.regfile_1.regOut[28] [6]),
    .R(rst_bF$buf25),
    .S(vdd)
);

FILL FILL_0__18823_ (
);

FILL FILL_0__18403_ (
);

OR2X2 _9669_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_631_)
);

OR2X2 _9249_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_411_)
);

FILL FILL370120x232180 (
);

FILL FILL_0__8924_ (
);

FILL FILL_0__8504_ (
);

FILL FILL_1__14389_ (
);

FILL FILL_1_BUFX2_insert1060 (
);

OR2X2 _13667_ (
    .A(_3151_),
    .B(_3148_),
    .Y(\datapath_1.mux_pcsrc.dout [10])
);

AND2X2 _13247_ (
    .A(_2791_),
    .B(_2233_),
    .Y(_2792_)
);

FILL FILL_1_BUFX2_insert1068 (
);

OR2X2 _17080_ (
    .A(_5994_),
    .B(_6009_),
    .Y(_6010_)
);

FILL FILL_0__9709_ (
);

FILL FILL271320x9880 (
);

FILL FILL_1__16535_ (
);

FILL FILL143640x34580 (
);

FILL FILL_0__15528_ (
);

AND2X2 _15813_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_4762_)
);

FILL FILL_0__15108_ (
);

FILL FILL_0__10663_ (
);

FILL FILL137560x172900 (
);

OR2X2 _18285_ (
    .A(_7182_),
    .B(_7196_),
    .Y(_7197_)
);

FILL FILL150480x167960 (
);

FILL FILL254600x4940 (
);

FILL FILL_0__9882_ (
);

FILL FILL_0__11448_ (
);

FILL FILL_0__9042_ (
);

OR2X2 _11733_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_1687_)
);

OR2X2 _11313_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_1467_)
);

FILL FILL_0__15281_ (
);

FILL FILL212040x192660 (
);

FILL FILL273600x4940 (
);

FILL FILL_1_BUFX2_insert680 (
);

AOI21X1 _12938_ (
    .A(_2164_),
    .B(_2161_),
    .C(_2501_),
    .Y(_2502_)
);

INVX1 _12518_ (
    .A(_2108_),
    .Y(_2109_)
);

FILL FILL_1_BUFX2_insert688 (
);

FILL FILL_0__16486_ (
);

AND2X2 _16771_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_5705_)
);

OR2X2 _16351_ (
    .A(_5290_),
    .B(_5291_),
    .Y(_5292_)
);

FILL FILL292600x4940 (
);

FILL FILL131480x113620 (
);

DFFSR _8693_ (
    .CLK(clk_bF$buf79),
    .D(_69_[11]),
    .Q(\datapath_1.regfile_1.regOut[2] [11]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL376960x44460 (
);

BUFX2 BUFX2_insert350 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf0 )
);

BUFX2 BUFX2_insert351 (
    .A(_3352_),
    .Y(_3352__bF$buf4)
);

BUFX2 BUFX2_insert352 (
    .A(_3352_),
    .Y(_3352__bF$buf3)
);

BUFX2 BUFX2_insert353 (
    .A(_3352_),
    .Y(_3352__bF$buf2)
);

BUFX2 BUFX2_insert354 (
    .A(_3352_),
    .Y(_3352__bF$buf1)
);

INVX1 _17976_ (
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_6893_)
);

FILL FILL471200x306280 (
);

AND2X2 _17556_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_6479_)
);

BUFX2 BUFX2_insert355 (
    .A(_3352_),
    .Y(_3352__bF$buf0)
);

BUFX2 BUFX2_insert356 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf4 )
);

AND2X2 _17136_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_6065_)
);

BUFX2 BUFX2_insert357 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf3 )
);

BUFX2 BUFX2_insert358 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf2 )
);

AND2X2 _12691_ (
    .A(_2253_),
    .B(_2255_),
    .Y(_2256_)
);

BUFX2 BUFX2_insert359 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf1 )
);

FILL FILL357200x330980 (
);

OR2X2 _12271_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .B(_1982__bF$buf3),
    .Y(_1966_)
);

FILL FILL249280x103740 (
);

OR2X2 _9898_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .B(_794__bF$buf0),
    .Y(_744_)
);

DFFSR _9478_ (
    .CLK(clk_bF$buf74),
    .D(_465_[22]),
    .Q(\datapath_1.regfile_1.regOut[8] [22]),
    .R(rst_bF$buf47),
    .S(vdd)
);

OR2X2 _9058_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .B(_332__bF$buf1),
    .Y(_324_)
);

FILL FILL_0__8733_ (
);

FILL FILL504640x24700 (
);

FILL FILL179360x108680 (
);

AND2X2 _13896_ (
    .A(_3330_),
    .B(_3329_),
    .Y(\datapath_1.alu_1.ALUInA [26])
);

OR2X2 _13476_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [19]),
    .Y(_3007_)
);

INVX1 _13056_ (
    .A(_2264_),
    .Y(_2613_)
);

FILL FILL236360x83980 (
);

FILL FILL_0__19417_ (
);

FILL FILL_0__14972_ (
);

FILL FILL_0__14552_ (
);

FILL FILL_0__14132_ (
);

FILL FILL_0__9938_ (
);

FILL FILL_0__9518_ (
);

FILL FILL105640x316160 (
);

FILL FILL_0__15757_ (
);

AND2X2 _15622_ (
    .A(_4223__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_4574_)
);

AND2X2 _15202_ (
    .A(_4141_),
    .B(_4128_),
    .Y(_4160_)
);

FILL FILL_0__10472_ (
);

FILL FILL_0__10052_ (
);

OR2X2 _18094_ (
    .A(_7007_),
    .B(_7008_),
    .Y(_7009_)
);

FILL FILL281960x197600 (
);

FILL FILL287280x271700 (
);

FILL FILL_0__19170_ (
);

FILL FILL_1__17549_ (
);

AND2X2 _16827_ (
    .A(_4217__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_5760_)
);

OR2X2 _16407_ (
    .A(_5343_),
    .B(_5346_),
    .Y(_5347_)
);

FILL FILL_0__9271_ (
);

OR2X2 _11962_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .B(_1850__bF$buf2),
    .Y(_1800_)
);

FILL FILL313120x266760 (
);

DFFSR _11542_ (
    .CLK(clk_bF$buf84),
    .D(_1521_[22]),
    .Q(\datapath_1.regfile_1.regOut[24] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

OR2X2 _11122_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .B(_1388__bF$buf0),
    .Y(_1380_)
);

INVX1 _19299_ (
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_8195_)
);

FILL FILL_0__17903_ (
);

FILL FILL467400x242060 (
);

OR2X2 _8749_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .B(_200__bF$buf2),
    .Y(_158_)
);

FILL FILL250040x44460 (
);

FILL FILL338960x74100 (
);

INVX1 _12747_ (
    .A(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2312_)
);

INVX2 _12327_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .Y(_2048_)
);

FILL FILL313880x251940 (
);

FILL FILL27360x237120 (
);

FILL FILL_0__13403_ (
);

FILL FILL213560x345800 (
);

OR2X2 _16580_ (
    .A(_5515_),
    .B(_5516_),
    .Y(_5517_)
);

FILL FILL_0__16295_ (
);

OR2X2 _16160_ (
    .A(_5100_),
    .B(_5103_),
    .Y(_5104_)
);

FILL FILL_1__9432_ (
);

FILL FILL367840x321100 (
);

FILL FILL_1__10330_ (
);

FILL FILL184680x14820 (
);

AND2X2 _17785_ (
    .A(_6289__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_6705_)
);

OR2X2 _17365_ (
    .A(_6288_),
    .B(_6290_),
    .Y(_6291_)
);

AND2X2 _12080_ (
    .A(_1858_),
    .B(_1857_),
    .Y(_1851_[3])
);

FILL FILL_0__18441_ (
);

FILL FILL_0__18021_ (
);

FILL FILL305520x281580 (
);

FILL FILL296400x177840 (
);

FILL FILL311600x222300 (
);

AND2X2 _9287_ (
    .A(_436_),
    .B(_435_),
    .Y(_399_[18])
);

FILL FILL164160x79040 (
);

OR2X2 _10813_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .B(_1256__bF$buf3),
    .Y(_1214_)
);

AND2X2 _13285_ (
    .A(_2824_),
    .B(_2827_),
    .Y(_2828_)
);

OR2X2 _19511_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_8376_)
);

FILL FILL209000x296400 (
);

FILL FILL_0__9747_ (
);

FILL FILL22040x88920 (
);

FILL FILL_1__16153_ (
);

FILL FILL_0__15986_ (
);

OR2X2 _15851_ (
    .A(_4798_),
    .B(_4799_),
    .Y(_4800_)
);

FILL FILL_0__15146_ (
);

OR2X2 _15431_ (
    .A(_4384_),
    .B(_4385_),
    .Y(_4386_)
);

DFFSR _15011_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[30]),
    .Q(\datapath_1.PCJump [30]),
    .R(rst_bF$buf18),
    .S(vdd)
);

FILL FILL_0__10281_ (
);

FILL FILL290320x118560 (
);

FILL FILL_1__12493_ (
);

AND2X2 _16636_ (
    .A(_4158__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_5572_)
);

OR2X2 _16216_ (
    .A(_5151_),
    .B(_5158_),
    .Y(_5159_)
);

FILL FILL_0__11486_ (
);

AND2X2 _11771_ (
    .A(_1712_),
    .B(_1711_),
    .Y(_1653_[29])
);

AND2X2 _11351_ (
    .A(_1492_),
    .B(_1491_),
    .Y(_1455_[18])
);

FILL FILL36480x355680 (
);

AND2X2 _8978_ (
    .A(_270_),
    .B(_269_),
    .Y(_267_[1])
);

DFFSR _8558_ (
    .CLK(clk_bF$buf59),
    .D(_3_[5]),
    .Q(\datapath_1.regfile_1.regOut[1] [5]),
    .R(rst_bF$buf106),
    .S(vdd)
);

FILL FILL102600x350740 (
);

FILL FILL275120x197600 (
);

AND2X2 _12976_ (
    .A(_2537_),
    .B(_2530_),
    .Y(_2538_)
);

NOR2X1 _12556_ (
    .A(_2107_),
    .B(_2105_),
    .Y(_2077_)
);

OR2X2 _12136_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .B(_1916__bF$buf3),
    .Y(_1896_)
);

FILL FILL_0__18917_ (
);

FILL FILL_0__13632_ (
);

FILL FILL_0__13212_ (
);

FILL FILL_1__9241_ (
);

FILL FILL_0__14837_ (
);

FILL FILL467400x24700 (
);

OR2X2 _14702_ (
    .A(vdd),
    .B(\datapath_1.a [25]),
    .Y(_3854_)
);

FILL FILL_0__14417_ (
);

BUFX2 BUFX2_insert730 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf3 )
);

BUFX2 BUFX2_insert731 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf2 )
);

BUFX2 BUFX2_insert732 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf1 )
);

BUFX2 BUFX2_insert733 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf0 )
);

BUFX2 BUFX2_insert734 (
    .A(_4183_),
    .Y(_4183__bF$buf4)
);

BUFX2 BUFX2_insert735 (
    .A(_4183_),
    .Y(_4183__bF$buf3)
);

AND2X2 _17594_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_6517_)
);

BUFX2 BUFX2_insert736 (
    .A(_4183_),
    .Y(_4183__bF$buf2)
);

OR2X2 _17174_ (
    .A(_6101_),
    .B(_6100_),
    .Y(_6102_)
);

BUFX2 BUFX2_insert737 (
    .A(_4183_),
    .Y(_4183__bF$buf1)
);

BUFX2 BUFX2_insert738 (
    .A(_4183_),
    .Y(_4183__bF$buf0)
);

FILL FILL503880x306280 (
);

BUFX2 BUFX2_insert739 (
    .A(_4239_),
    .Y(_4239__bF$buf4)
);

FILL FILL20520x350740 (
);

FILL FILL_0__18670_ (
);

FILL FILL_0__18250_ (
);

FILL FILL324520x261820 (
);

DFFSR _9096_ (
    .CLK(clk_bF$buf36),
    .D(_267_[27]),
    .Q(\datapath_1.regfile_1.regOut[5] [27]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL_1__11764_ (
);

FILL FILL332880x4940 (
);

OR2X2 _15907_ (
    .A(_4854_),
    .B(_4853_),
    .Y(_4855_)
);

FILL FILL_0__10337_ (
);

DFFSR _10622_ (
    .CLK(clk_bF$buf68),
    .D(_1059_[5]),
    .Q(\datapath_1.regfile_1.regOut[17] [5]),
    .R(rst_bF$buf40),
    .S(vdd)
);

AND2X2 _10202_ (
    .A(_906_),
    .B(_905_),
    .Y(_861_[22])
);

INVX1 _18799_ (
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_7703_)
);

OR2X2 _18379_ (
    .A(_7288_),
    .B(_7289_),
    .Y(_7290_)
);

FILL FILL83600x0 (
);

AND2X2 _13094_ (
    .A(_2647_),
    .B(_2648_),
    .Y(_2649_)
);

FILL FILL444600x98800 (
);

FILL FILL_0__19455_ (
);

FILL FILL_0__19035_ (
);

AND2X2 _19320_ (
    .A(_6262__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_8216_)
);

FILL FILL_0__14590_ (
);

FILL FILL_0__14170_ (
);

FILL FILL_1__12129_ (
);

FILL FILL274360x74100 (
);

FILL FILL351880x4940 (
);

FILL FILL_0__9556_ (
);

OR2X2 _11827_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .B(_1784__bF$buf1),
    .Y(_1730_)
);

DFFSR _11407_ (
    .CLK(clk_bF$buf0),
    .D(_1455_[16]),
    .Q(\datapath_1.regfile_1.regOut[23] [16]),
    .R(rst_bF$buf95),
    .S(vdd)
);

AND2X2 _14299_ (
    .A(_3645_),
    .B(_3644_),
    .Y(_3606_[19])
);

FILL FILL_0__12903_ (
);

FILL FILL_0__15795_ (
);

FILL FILL_0__15375_ (
);

AND2X2 _15660_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_4612_)
);

AND2X2 _15240_ (
    .A(_4197__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_4198_)
);

FILL FILL_0__10090_ (
);

AND2X2 _16865_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_5798_)
);

OR2X2 _16445_ (
    .A(_5382_),
    .B(_5383_),
    .Y(_5384_)
);

OR2X2 _16025_ (
    .A(_4955_),
    .B(_4970_),
    .Y(_4971_)
);

OR2X2 _11580_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_1605_)
);

DFFSR _11160_ (
    .CLK(clk_bF$buf68),
    .D(_1323_[27]),
    .Q(\datapath_1.regfile_1.regOut[21] [27]),
    .R(rst_bF$buf40),
    .S(vdd)
);

FILL FILL23560x29640 (
);

FILL FILL_0__17941_ (
);

FILL FILL_0__17521_ (
);

OR2X2 _8787_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_183_)
);

FILL FILL424080x19760 (
);

FILL FILL298680x276640 (
);

FILL FILL_1__13087_ (
);

AND2X2 _12785_ (
    .A(_2338_),
    .B(_2349_),
    .Y(_2350_)
);

AND2X2 _12365_ (
    .A(_2008_),
    .B(_2007_),
    .Y(_1983_[12])
);

FILL FILL_1__19313_ (
);

FILL FILL_0__18306_ (
);

FILL FILL_0__13861_ (
);

FILL FILL_0__13021_ (
);

FILL FILL_1__9050_ (
);

FILL FILL66120x207480 (
);

FILL FILL256120x370500 (
);

FILL FILL_1__15653_ (
);

FILL FILL47120x365560 (
);

FILL FILL_0__14646_ (
);

OR2X2 _14931_ (
    .A(\datapath_1.mux_pcsrc.dout [15]),
    .B(_4001__bF$buf3),
    .Y(_3967_)
);

FILL FILL_0__14226_ (
);

OR2X2 _14511_ (
    .A(memoryOutData[4]),
    .B(_3803__bF$buf2),
    .Y(_3747_)
);

FILL FILL96520x163020 (
);

FILL FILL210520x311220 (
);

FILL FILL_1__16018_ (
);

FILL FILL368600x286520 (
);

FILL FILL_1__11573_ (
);

AND2X2 _15716_ (
    .A(_4208__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_4667_)
);

FILL FILL_0__10986_ (
);

OR2X2 _10851_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_1239_)
);

OR2X2 _10431_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_1019_)
);

FILL FILL_0__10146_ (
);

OR2X2 _10011_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_799_)
);

OR2X2 _18188_ (
    .A(_7069_),
    .B(_7101_),
    .Y(_7102_)
);

FILL FILL_0__19264_ (
);

FILL FILL_1__12778_ (
);

FILL FILL104880x128440 (
);

FILL FILL_0__9785_ (
);

FILL FILL_0__9365_ (
);

AND2X2 _11636_ (
    .A(_1642_),
    .B(_1641_),
    .Y(_1587_[27])
);

AND2X2 _11216_ (
    .A(_1422_),
    .B(_1421_),
    .Y(_1389_[16])
);

FILL FILL250040x311220 (
);

FILL FILL_0__12712_ (
);

FILL FILL_1__8741_ (
);

FILL FILL108680x370500 (
);

FILL FILL462840x133380 (
);

FILL FILL504640x261820 (
);

AND2X2 _16674_ (
    .A(_4167__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_5610_)
);

AND2X2 _16254_ (
    .A(_4189__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_5196_)
);

FILL FILL62320x237120 (
);

FILL FILL385320x311220 (
);

OR2X2 _8596_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .B(_134__bF$buf4),
    .Y(_76_)
);

FILL FILL371640x9880 (
);

OR2X2 _17879_ (
    .A(_6796_),
    .B(_6795_),
    .Y(_6797_)
);

OR2X2 _17459_ (
    .A(_6382_),
    .B(_6383_),
    .Y(_6384_)
);

OR2X2 _17039_ (
    .A(_5968_),
    .B(_5967_),
    .Y(_5969_)
);

NAND2X1 _12594_ (
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2159_)
);

DFFSR _12174_ (
    .CLK(clk_bF$buf72),
    .D(_1851_[9]),
    .Q(\datapath_1.regfile_1.regOut[29] [9]),
    .R(rst_bF$buf2),
    .S(vdd)
);

FILL FILL380000x98800 (
);

FILL FILL_0__18955_ (
);

OR2X2 _18820_ (
    .A(_7720_),
    .B(_7723_),
    .Y(_7724_)
);

FILL FILL_0__18535_ (
);

FILL FILL_0__18115_ (
);

OR2X2 _18400_ (
    .A(_7302_),
    .B(_7309_),
    .Y(_7310_)
);

FILL FILL_0__13250_ (
);

FILL FILL_0__8636_ (
);

OR2X2 _10907_ (
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .Y(_1321_)
);

FILL FILL119320x108680 (
);

FILL FILL190000x0 (
);

OR2X2 _13799_ (
    .A(_3264_),
    .B(_3263_),
    .Y(_3265_)
);

AND2X2 _13379_ (
    .A(_2916_),
    .B(_2914_),
    .Y(_2917_)
);

FILL FILL_1__15042_ (
);

DFFSR _14740_ (
    .CLK(clk_bF$buf40),
    .D(_3804_[17]),
    .Q(\datapath_1.a [17]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL_0__14035_ (
);

AND2X2 _14320_ (
    .A(_3659_),
    .B(_3658_),
    .Y(_3606_[26])
);

FILL FILL424080x143260 (
);

FILL FILL223440x350740 (
);

FILL FILL309320x365560 (
);

FILL FILL_1__11382_ (
);

OR2X2 _15945_ (
    .A(_4891_),
    .B(_4884_),
    .Y(_4892_)
);

AND2X2 _15525_ (
    .A(_4197__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_4479_)
);

NAND3X1 _15105_ (
    .A(_4013_),
    .B(_4002_),
    .C(_4017_),
    .Y(_4086_)
);

FILL FILL_0__10795_ (
);

OR2X2 _10660_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .B(_1190__bF$buf2),
    .Y(_1132_)
);

DFFSR _10240_ (
    .CLK(clk_bF$buf33),
    .D(_861_[10]),
    .Q(\datapath_1.regfile_1.regOut[14] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

FILL FILL153520x355680 (
);

FILL FILL_0__16601_ (
);

FILL FILL326800x375440 (
);

FILL FILL_0__19493_ (
);

FILL FILL218880x148200 (
);

FILL FILL240160x266760 (
);

FILL FILL54720x118560 (
);

FILL FILL_1__18813_ (
);

OR2X2 _11865_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_1755_)
);

FILL FILL_0__9174_ (
);

OR2X2 _11445_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_1535_)
);

DFFSR _11025_ (
    .CLK(clk_bF$buf47),
    .D(_1257_[21]),
    .Q(\datapath_1.regfile_1.regOut[20] [21]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL_0__12521_ (
);

FILL FILL_0__12101_ (
);

FILL FILL339720x187720 (
);

FILL FILL476520x247000 (
);

FILL FILL_0__13726_ (
);

FILL FILL_0_BUFX2_insert1070 (
);

FILL FILL_0_BUFX2_insert1072 (
);

OR2X2 _16483_ (
    .A(_5421_),
    .B(_5420_),
    .Y(_5422_)
);

FILL FILL_0__16198_ (
);

AND2X2 _16063_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_5008_)
);

FILL FILL_0_BUFX2_insert1074 (
);

FILL FILL_0_BUFX2_insert1075 (
);

FILL FILL_0_BUFX2_insert1076 (
);

FILL FILL_0_BUFX2_insert1077 (
);

FILL FILL_0_BUFX2_insert1078 (
);

FILL FILL75240x276640 (
);

FILL FILL160360x242060 (
);

FILL FILL_1__15518_ (
);

FILL FILL133760x74100 (
);

FILL FILL150480x24700 (
);

AND2X2 _17688_ (
    .A(_6247__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_6609_)
);

AND2X2 _17268_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_6195_)
);

FILL FILL_0__18764_ (
);

FILL FILL_0__18344_ (
);

FILL FILL342000x251940 (
);

FILL FILL_0__8865_ (
);

FILL FILL_0__8445_ (
);

OR2X2 _10716_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_1169_)
);

NAND3X1 _13188_ (
    .A(_2379__bF$buf1),
    .B(\datapath_1.alu_1.ALUInB [15]),
    .C(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2737_)
);

FILL FILL_1__15271_ (
);

AND2X2 _19414_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_8309_)
);

FILL FILL_0__19129_ (
);

FILL FILL11400x98800 (
);

FILL FILL505400x0 (
);

FILL FILL154280x24700 (
);

FILL FILL_1__16476_ (
);

FILL FILL_1__11191_ (
);

AND2X2 _15754_ (
    .A(_4214__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_4704_)
);

FILL FILL_0__15469_ (
);

FILL FILL_0__15049_ (
);

OR2X2 _15334_ (
    .A(_4290_),
    .B(_4289_),
    .Y(_4291_)
);

FILL FILL50160x375440 (
);

FILL FILL_0__10184_ (
);

FILL FILL_0__16410_ (
);

FILL FILL354160x286520 (
);

AND2X2 _16959_ (
    .A(_4146__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_5890_)
);

AND2X2 _16539_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_5477_)
);

OR2X2 _16119_ (
    .A(_5056_),
    .B(_5063_),
    .Y(_5064_)
);

FILL FILL_0__11389_ (
);

DFFSR _11674_ (
    .CLK(clk_bF$buf60),
    .D(_1587_[25]),
    .Q(\datapath_1.regfile_1.regOut[25] [25]),
    .R(rst_bF$buf101),
    .S(vdd)
);

OR2X2 _11254_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_1454__bF$buf4),
    .Y(_1448_)
);

FILL FILL6840x167960 (
);

FILL FILL52440x74100 (
);

FILL FILL_0__17615_ (
);

AND2X2 _17900_ (
    .A(_6289__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_6818_)
);

FILL FILL_0__12750_ (
);

FILL FILL_0__12330_ (
);

OR2X2 _9822_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_713_)
);

OR2X2 _9402_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_493_)
);

FILL FILL452200x163020 (
);

OR2X2 _12879_ (
    .A(_2443_),
    .B(_2419_),
    .Y(_2444_)
);

NAND2X1 _12459_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2053_)
);

DFFSR _12039_ (
    .CLK(clk_bF$buf46),
    .D(_1785_[3]),
    .Q(\datapath_1.regfile_1.regOut[28] [3]),
    .R(rst_bF$buf97),
    .S(vdd)
);

FILL FILL278920x232180 (
);

OR2X2 _13820_ (
    .A(\datapath_1.a [1]),
    .B(_3342__bF$buf1),
    .Y(_3280_)
);

FILL FILL_0__13115_ (
);

XOR2X1 _13400_ (
    .A(_2392_),
    .B(_2181_),
    .Y(_2936_)
);

AND2X2 _16292_ (
    .A(_4146__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_5234_)
);

FILL FILL329080x291460 (
);

FILL FILL178600x326040 (
);

FILL FILL96520x24700 (
);

FILL FILL_1__9144_ (
);

FILL FILL164920x350740 (
);

FILL FILL_1__10462_ (
);

DFFSR _14605_ (
    .CLK(clk_bF$buf23),
    .D(_3738_[11]),
    .Q(\datapath_1.PCJump [13]),
    .R(rst_bF$buf33),
    .S(vdd)
);

FILL FILL372400x93860 (
);

AND2X2 _17497_ (
    .A(_6236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_6421_)
);

FILL FILL280440x0 (
);

OR2X2 _17077_ (
    .A(_6005_),
    .B(_6006_),
    .Y(_6007_)
);

FILL FILL_0__18993_ (
);

FILL FILL486400x182780 (
);

FILL FILL_0__18573_ (
);

FILL FILL346560x167960 (
);

OR2X2 _10945_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_1322__bF$buf1),
    .Y(_1282_)
);

OR2X2 _10525_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .B(_1124__bF$buf0),
    .Y(_1062_)
);

DFFSR _10105_ (
    .CLK(clk_bF$buf73),
    .D(_795_[4]),
    .Q(\datapath_1.regfile_1.regOut[13] [4]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL105640x202540 (
);

FILL FILL_0__11601_ (
);

FILL FILL46360x177840 (
);

FILL FILL_0__19358_ (
);

AND2X2 _19223_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_8121_)
);

FILL FILL_0__14073_ (
);

FILL FILL_0__9879_ (
);

FILL FILL386840x261820 (
);

FILL FILL203680x182780 (
);

OR2X2 _15983_ (
    .A(_4926_),
    .B(_4929_),
    .Y(_4930_)
);

FILL FILL_0__15698_ (
);

FILL FILL_0__15278_ (
);

AND2X2 _15563_ (
    .A(_4197__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_4516_)
);

NOR2X1 _15143_ (
    .A(_4110_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.regfile_1.regEn [22])
);

FILL FILL199880x335920 (
);

FILL FILL340480x108680 (
);

OR2X2 _16768_ (
    .A(_5701_),
    .B(_5700_),
    .Y(_5702_)
);

OR2X2 _16348_ (
    .A(_5287_),
    .B(_5288_),
    .Y(_5289_)
);

FILL FILL380000x217360 (
);

FILL FILL143640x370500 (
);

AND2X2 _11483_ (
    .A(_1560_),
    .B(_1559_),
    .Y(_1521_[19])
);

FILL FILL_1__18431_ (
);

FILL FILL_0__11198_ (
);

AND2X2 _11063_ (
    .A(_1340_),
    .B(_1339_),
    .Y(_1323_[8])
);

FILL FILL_0__17424_ (
);

FILL FILL_0__17004_ (
);

FILL FILL38760x192660 (
);

OR2X2 _9631_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .B(_662__bF$buf2),
    .Y(_606_)
);

DFFSR _9211_ (
    .CLK(clk_bF$buf52),
    .D(_333_[13]),
    .Q(\datapath_1.regfile_1.regOut[6] [13]),
    .R(rst_bF$buf90),
    .S(vdd)
);

FILL FILL21280x276640 (
);

NAND3X1 _12688_ (
    .A(_2211_),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .C(_2252_),
    .Y(_2253_)
);

OR2X2 _12268_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .B(_1982__bF$buf4),
    .Y(_1964_)
);

FILL FILL_0__18629_ (
);

AND2X2 _18914_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_7816_)
);

FILL FILL_0__18209_ (
);

FILL FILL_0__13764_ (
);

FILL FILL_0__13344_ (
);

FILL FILL348080x271700 (
);

FILL FILL505400x158080 (
);

FILL FILL224200x103740 (
);

FILL FILL_1__15136_ (
);

FILL FILL_1__10271_ (
);

FILL FILL278160x276640 (
);

OR2X2 _14834_ (
    .A(vdd),
    .B(_2_[26]),
    .Y(_3922_)
);

FILL FILL_0__14549_ (
);

OR2X2 _14414_ (
    .A(vdd),
    .B(\datapath_1.Data [15]),
    .Y(_3702_)
);

FILL FILL162640x34580 (
);

FILL FILL_0__15910_ (
);

FILL FILL372400x232180 (
);

FILL FILL_0__18382_ (
);

FILL FILL269800x19760 (
);

AND2X2 _15619_ (
    .A(_4197__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_4571_)
);

FILL FILL_0__8483_ (
);

DFFSR _10754_ (
    .CLK(clk_bF$buf63),
    .D(_1125_[8]),
    .Q(\datapath_1.regfile_1.regOut[18] [8]),
    .R(rst_bF$buf58),
    .S(vdd)
);

FILL FILL_0__10469_ (
);

FILL FILL_0__10049_ (
);

AND2X2 _10334_ (
    .A(_974_),
    .B(_973_),
    .Y(_927_[23])
);

FILL FILL72200x242060 (
);

FILL FILL376200x153140 (
);

OR2X2 _19452_ (
    .A(gnd),
    .B(_8385__bF$buf1),
    .Y(_8337_)
);

OR2X2 _19032_ (
    .A(_7932_),
    .B(_7916_),
    .Y(_7933_)
);

OR2X2 _8902_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .B(_266__bF$buf1),
    .Y(_240_)
);

FILL FILL_0__9688_ (
);

FILL FILL185440x306280 (
);

FILL FILL_0__9268_ (
);

OR2X2 _11959_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_1850__bF$buf2),
    .Y(_1798_)
);

DFFSR _11539_ (
    .CLK(clk_bF$buf80),
    .D(_1521_[19]),
    .Q(\datapath_1.regfile_1.regOut[24] [19]),
    .R(rst_bF$buf76),
    .S(vdd)
);

FILL FILL327560x340860 (
);

OR2X2 _11119_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .B(_1388__bF$buf3),
    .Y(_1378_)
);

FILL FILL_1__13622_ (
);

FILL FILL_1_BUFX2_insert300 (
);

OR2X2 _12900_ (
    .A(_2452_),
    .B(_2464_),
    .Y(_2465_)
);

FILL FILL_0__12615_ (
);

FILL FILL_1__16094_ (
);

FILL FILL_1_BUFX2_insert309 (
);

AND2X2 _15792_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_4742_)
);

FILL FILL_0__15087_ (
);

OR2X2 _15372_ (
    .A(_4327_),
    .B(_4326_),
    .Y(_4328_)
);

FILL FILL_1__14827_ (
);

FILL FILL411920x49400 (
);

AND2X2 _16997_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_5928_)
);

OR2X2 _16577_ (
    .A(_5510_),
    .B(_5513_),
    .Y(_5514_)
);

AND2X2 _16157_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_5101_)
);

DFFSR _11292_ (
    .CLK(clk_bF$buf54),
    .D(_1389_[30]),
    .Q(\datapath_1.regfile_1.regOut[22] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL_0__17653_ (
);

FILL FILL_0__17233_ (
);

OR2X2 _8499_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_31_)
);

FILL FILL183920x0 (
);

DFFSR _9860_ (
    .CLK(clk_bF$buf109),
    .D(_663_[17]),
    .Q(\datapath_1.regfile_1.regOut[11] [17]),
    .R(rst_bF$buf64),
    .S(vdd)
);

AND2X2 _9440_ (
    .A(_518_),
    .B(_517_),
    .Y(_465_[26])
);

FILL FILL57760x172900 (
);

AND2X2 _9020_ (
    .A(_298_),
    .B(_297_),
    .Y(_267_[15])
);

FILL FILL205200x167960 (
);

NAND2X1 _12497_ (
    .A(_2094_),
    .B(_2098_),
    .Y(ALUSrcA)
);

AND2X2 _12077_ (
    .A(_1856_),
    .B(_1855_),
    .Y(_1851_[2])
);

FILL FILL_1__14580_ (
);

FILL FILL_0__18858_ (
);

AND2X2 _18723_ (
    .A(_6221__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_7628_)
);

FILL FILL_0__18438_ (
);

AND2X2 _18303_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_7215_)
);

FILL FILL_0__13993_ (
);

FILL FILL_0__13573_ (
);

FILL FILL_0__13153_ (
);

FILL FILL293360x335920 (
);

FILL FILL133760x113620 (
);

FILL FILL128440x247000 (
);

FILL FILL_0__8539_ (
);

FILL FILL_1__9182_ (
);

OR2X2 _19508_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_8374_)
);

FILL FILL_0__14778_ (
);

OR2X2 _14643_ (
    .A(\datapath_1.rd1 [5]),
    .B(_3869__bF$buf3),
    .Y(_3815_)
);

FILL FILL306280x360620 (
);

AND2X2 _14223_ (
    .A(_3593_),
    .B(_3592_),
    .Y(\datapath_1.mux_wd3.dout [26])
);

FILL FILL351880x103740 (
);

FILL FILL128440x64220 (
);

FILL FILL437760x118560 (
);

OR2X2 _15848_ (
    .A(_4796_),
    .B(_4789_),
    .Y(_4797_)
);

OR2X2 _15428_ (
    .A(_4382_),
    .B(_4381_),
    .Y(_4383_)
);

DFFSR _15008_ (
    .CLK(clk_bF$buf92),
    .D(_3936_[27]),
    .Q(\datapath_1.mux_iord.din0 [27]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL_1__17931_ (
);

OR2X2 _10983_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_1307_)
);

OR2X2 _10563_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_1087_)
);

FILL FILL_0__10278_ (
);

OR2X2 _10143_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_867_)
);

FILL FILL_0__16504_ (
);

FILL FILL389120x192660 (
);

FILL FILL_0__19396_ (
);

AND2X2 _19261_ (
    .A(_6282__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_8158_)
);

FILL FILL38760x9880 (
);

DFFSR _8711_ (
    .CLK(clk_bF$buf30),
    .D(_69_[29]),
    .Q(\datapath_1.regfile_1.regOut[2] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

FILL FILL_0__9497_ (
);

AND2X2 _11768_ (
    .A(_1710_),
    .B(_1709_),
    .Y(_1653_[28])
);

AND2X2 _11348_ (
    .A(_1490_),
    .B(_1489_),
    .Y(_1455_[17])
);

FILL FILL122360x88920 (
);

FILL FILL504640x98800 (
);

FILL FILL_1__13011_ (
);

FILL FILL_0__17709_ (
);

FILL FILL_0__12844_ (
);

FILL FILL69920x93860 (
);

FILL FILL_0__12004_ (
);

AND2X2 _15181_ (
    .A(_4138_),
    .B(\datapath_1.PCJump [20]),
    .Y(_4139_)
);

OR2X2 _9916_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .B(_794__bF$buf1),
    .Y(_756_)
);

FILL FILL_1__8873_ (
);

FILL FILL289560x271700 (
);

FILL FILL_1__14636_ (
);

AND2X2 _13914_ (
    .A(_3344__bF$buf2),
    .B(gnd),
    .Y(_3345_)
);

FILL FILL_0__13629_ (
);

FILL FILL_0__13209_ (
);

AND2X2 _16386_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_5326_)
);

FILL FILL149720x88920 (
);

FILL FILL412680x217360 (
);

FILL FILL_0__17882_ (
);

FILL FILL_0__17462_ (
);

FILL FILL_0__17042_ (
);

FILL FILL338200x350740 (
);

FILL FILL383040x133380 (
);

FILL FILL233320x172900 (
);

FILL FILL319200x187720 (
);

FILL FILL183160x79040 (
);

FILL FILL_1__19254_ (
);

FILL FILL_0__10910_ (
);

AND2X2 _18952_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [24]),
    .Y(_7854_)
);

AND2X2 _18532_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_7440_)
);

OR2X2 _18112_ (
    .A(_7025_),
    .B(_7026_),
    .Y(_7027_)
);

FILL FILL_0__8768_ (
);

DFFSR _10619_ (
    .CLK(clk_bF$buf18),
    .D(_1059_[2]),
    .Q(\datapath_1.regfile_1.regOut[17] [2]),
    .R(rst_bF$buf107),
    .S(vdd)
);

FILL FILL_1__15594_ (
);

FILL FILL319960x59280 (
);

AND2X2 _19317_ (
    .A(_6259__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_8213_)
);

DFFSR _14872_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[20]),
    .Q(_2_[20]),
    .R(rst_bF$buf61),
    .S(vdd)
);

FILL FILL_0__14587_ (
);

FILL FILL_0__14167_ (
);

AND2X2 _14452_ (
    .A(_3727_),
    .B(_3726_),
    .Y(_3672_[27])
);

OR2X2 _14032_ (
    .A(_3445_),
    .B(_3446_),
    .Y(_3447_)
);

FILL FILL378480x118560 (
);

FILL FILL465880x123500 (
);

FILL FILL307800x281580 (
);

FILL FILL_1__13907_ (
);

FILL FILL252320x158080 (
);

FILL FILL505400x311220 (
);

FILL FILL313120x128440 (
);

AND2X2 _15657_ (
    .A(_4228__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_4609_)
);

NOR3X1 _15237_ (
    .A(_4150_),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .C(_4153_),
    .Y(_4195_)
);

OR2X2 _10792_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .B(_1256__bF$buf4),
    .Y(_1200_)
);

DFFSR _10372_ (
    .CLK(clk_bF$buf61),
    .D(_927_[13]),
    .Q(\datapath_1.regfile_1.regOut[15] [13]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL59280x286520 (
);

FILL FILL_0__16733_ (
);

FILL FILL155800x192660 (
);

OR2X2 _19490_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [21]),
    .Y(_8362_)
);

AND2X2 _19070_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_7970_)
);

DFFSR _8940_ (
    .CLK(clk_bF$buf35),
    .D(_201_[0]),
    .Q(\datapath_1.regfile_1.regOut[4] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

OR2X2 _8520_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_45_)
);

OR2X2 _11997_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_1823_)
);

OR2X2 _11577_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_1603_)
);

FILL FILL_1__18105_ (
);

DFFSR _11157_ (
    .CLK(clk_bF$buf97),
    .D(_1323_[24]),
    .Q(\datapath_1.regfile_1.regOut[21] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL_1__13660_ (
);

FILL FILL_0__17938_ (
);

OR2X2 _17803_ (
    .A(_6721_),
    .B(_6720_),
    .Y(_6722_)
);

FILL FILL_0__12233_ (
);

FILL FILL142120x197600 (
);

FILL FILL167200x49400 (
);

DFFSR _9725_ (
    .CLK(clk_bF$buf95),
    .D(_597_[11]),
    .Q(\datapath_1.regfile_1.regOut[10] [11]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL344280x326040 (
);

AND2X2 _9305_ (
    .A(_448_),
    .B(_447_),
    .Y(_399_[24])
);

FILL FILL56240x182780 (
);

FILL FILL_0__13858_ (
);

FILL FILL_0__13438_ (
);

OR2X2 _13723_ (
    .A(_3199_),
    .B(_3196_),
    .Y(\datapath_1.mux_pcsrc.dout [18])
);

OR2X2 _13303_ (
    .A(_2387__bF$buf2),
    .B(_2844_),
    .Y(_2845_)
);

FILL FILL_0__13018_ (
);

AND2X2 _16195_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_5138_)
);

FILL FILL38760x355680 (
);

FILL FILL_1__9887_ (
);

FILL FILL9880x153140 (
);

FILL FILL123880x29640 (
);

FILL FILL_0__17691_ (
);

FILL FILL369360x0 (
);

OR2X2 _14928_ (
    .A(\datapath_1.mux_pcsrc.dout [14]),
    .B(_4001__bF$buf0),
    .Y(_3965_)
);

OR2X2 _14508_ (
    .A(memoryOutData[3]),
    .B(_3803__bF$buf3),
    .Y(_3745_)
);

FILL FILL186960x256880 (
);

FILL FILL104120x256880 (
);

AND2X2 _18761_ (
    .A(_6289__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_7666_)
);

FILL FILL_0__18476_ (
);

OR2X2 _18341_ (
    .A(_7248_),
    .B(_7251_),
    .Y(_7252_)
);

FILL FILL_0__18056_ (
);

FILL FILL_0__13191_ (
);

FILL FILL121600x266760 (
);

FILL FILL_0__8997_ (
);

OR2X2 _10848_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_1237_)
);

OR2X2 _10428_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_1017_)
);

OR2X2 _10008_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_797_)
);

FILL FILL_0__11504_ (
);

FILL FILL127680x29640 (
);

DFFSR _19546_ (
    .CLK(clk_bF$buf84),
    .D(_8320_[23]),
    .Q(\datapath_1.regfile_1.regOut[0] [23]),
    .R(rst_bF$buf47),
    .S(vdd)
);

OR2X2 _19126_ (
    .A(_8024_),
    .B(_8023_),
    .Y(_8025_)
);

OR2X2 _14681_ (
    .A(vdd),
    .B(\datapath_1.a [18]),
    .Y(_3840_)
);

FILL FILL_0__14396_ (
);

OR2X2 _14261_ (
    .A(vdd),
    .B(ALUOut[7]),
    .Y(_3620_)
);

FILL FILL_0__12709_ (
);

FILL FILL326040x167960 (
);

AND2X2 _15886_ (
    .A(_4172__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_4834_)
);

AND2X2 _15466_ (
    .A(_4167__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_4421_)
);

NAND3X1 _15046_ (
    .A(_4031_),
    .B(_4017_),
    .C(_4012_),
    .Y(_4035_)
);

AND2X2 _10181_ (
    .A(_892_),
    .B(_891_),
    .Y(_861_[15])
);

FILL FILL_0__16542_ (
);

FILL FILL_0__16122_ (
);

FILL FILL76000x326040 (
);

FILL FILL279680x158080 (
);

FILL FILL114760x83980 (
);

FILL FILL_1__18754_ (
);

OR2X2 _11386_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .B(_1520__bF$buf3),
    .Y(_1516_)
);

FILL FILL_0__17747_ (
);

OR2X2 _17612_ (
    .A(_6533_),
    .B(_6530_),
    .Y(_6534_)
);

FILL FILL_0__17327_ (
);

FILL FILL_0__12882_ (
);

FILL FILL_0__12462_ (
);

FILL FILL338960x296400 (
);

OR2X2 _9954_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_781_)
);

FILL FILL278920x59280 (
);

OR2X2 _9534_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_561_)
);

OR2X2 _9114_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[6] [4]),
    .Y(_341_)
);

FILL FILL_1__19119_ (
);

AND2X2 _18817_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_7721_)
);

FILL FILL_0_BUFX2_insert340 (
);

FILL FILL231800x29640 (
);

FILL FILL_0_BUFX2_insert341 (
);

FILL FILL_0_BUFX2_insert342 (
);

FILL FILL_0_BUFX2_insert343 (
);

OR2X2 _13952_ (
    .A(_3378_),
    .B(_3375_),
    .Y(\datapath_1.alu_1.ALUInB [4])
);

FILL FILL_0__13667_ (
);

OR2X2 _13532_ (
    .A(ALUOut[14]),
    .B(_3079__bF$buf2),
    .Y(_3043_)
);

FILL FILL_0_BUFX2_insert345 (
);

INVX1 _13112_ (
    .A(_2284_),
    .Y(_2665_)
);

FILL FILL_0_BUFX2_insert347 (
);

FILL FILL_0_BUFX2_insert349 (
);

FILL FILL193040x9880 (
);

FILL FILL89680x123500 (
);

FILL FILL318440x182780 (
);

FILL FILL_1__9276_ (
);

FILL FILL_0__17080_ (
);

FILL FILL_1__15459_ (
);

FILL FILL_1__10594_ (
);

DFFSR _14737_ (
    .CLK(clk_bF$buf38),
    .D(_3804_[14]),
    .Q(\datapath_1.a [14]),
    .R(rst_bF$buf15),
    .S(vdd)
);

AND2X2 _14317_ (
    .A(_3657_),
    .B(_3656_),
    .Y(_3606_[25])
);

FILL FILL_1__16400_ (
);

OR2X2 _18990_ (
    .A(_7887_),
    .B(_7890_),
    .Y(_7891_)
);

AND2X2 _18570_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_7478_)
);

AND2X2 _18150_ (
    .A(_6315__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_7064_)
);

FILL FILL68400x207480 (
);

FILL FILL258400x370500 (
);

OR2X2 _10657_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .B(_1190__bF$buf4),
    .Y(_1130_)
);

DFFSR _10237_ (
    .CLK(clk_bF$buf29),
    .D(_861_[7]),
    .Q(\datapath_1.regfile_1.regOut[14] [7]),
    .R(rst_bF$buf21),
    .S(vdd)
);

FILL FILL_1__12740_ (
);

FILL FILL49400x365560 (
);

FILL FILL_0__11733_ (
);

FILL FILL_0__11313_ (
);

OR2X2 _19355_ (
    .A(_8247_),
    .B(_8250_),
    .Y(_8251_)
);

DFFSR _14490_ (
    .CLK(clk_bF$buf78),
    .D(_3672_[25]),
    .Q(\datapath_1.Data [25]),
    .R(rst_bF$buf26),
    .S(vdd)
);

OR2X2 _14070_ (
    .A(_3479_),
    .B(_3478_),
    .Y(_3480_)
);

OR2X2 _8805_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_195_)
);

FILL FILL125400x306280 (
);

FILL FILL212800x311220 (
);

FILL FILL294880x217360 (
);

FILL FILL_0__12938_ (
);

AND2X2 _12803_ (
    .A(_2366_),
    .B(_2367_),
    .Y(_2368_)
);

OR2X2 _15695_ (
    .A(_4644_),
    .B(_4645_),
    .Y(_4646_)
);

OR2X2 _15275_ (
    .A(_4227_),
    .B(_4232_),
    .Y(_4233_)
);

FILL FILL152000x59280 (
);

FILL FILL_1__8547_ (
);

FILL FILL_0__16771_ (
);

FILL FILL_0__16351_ (
);

FILL FILL252320x311220 (
);

AND2X2 _11195_ (
    .A(_1408_),
    .B(_1407_),
    .Y(_1389_[9])
);

FILL FILL_0__17976_ (
);

FILL FILL_0__17556_ (
);

OR2X2 _17841_ (
    .A(_6759_),
    .B(_6758_),
    .Y(_6760_)
);

AND2X2 _17421_ (
    .A(_6312__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_6346_)
);

AND2X2 _17001_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_5932_)
);

FILL FILL_0__12691_ (
);

FILL FILL505400x4940 (
);

OR2X2 _9763_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .B(_728__bF$buf2),
    .Y(_674_)
);

DFFSR _9343_ (
    .CLK(clk_bF$buf5),
    .D(_399_[16]),
    .Q(\datapath_1.regfile_1.regOut[7] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

FILL FILL10640x167960 (
);

FILL FILL_1__14063_ (
);

OR2X2 _18626_ (
    .A(_7525_),
    .B(_7532_),
    .Y(_7533_)
);

AND2X2 _18206_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_7119_)
);

OR2X2 _13761_ (
    .A(_3230_),
    .B(_3231_),
    .Y(_3232_)
);

FILL FILL_0__13056_ (
);

NOR2X1 _13341_ (
    .A(_2871_),
    .B(_2498_),
    .Y(_2881_)
);

FILL FILL64600x237120 (
);

FILL FILL387600x311220 (
);

FILL FILL3800x247000 (
);

FILL FILL_0__9803_ (
);

FILL FILL368600x148200 (
);

FILL FILL_1__15688_ (
);

FILL FILL349600x0 (
);

OR2X2 _14966_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [27]),
    .Y(_3990_)
);

OR2X2 _14546_ (
    .A(IRWrite_bF$buf4),
    .B(\datapath_1.PCJump [18]),
    .Y(_3770_)
);

OR2X2 _14126_ (
    .A(_3527_),
    .B(_3526_),
    .Y(_3528_)
);

FILL FILL_0__15622_ (
);

FILL FILL_0__15202_ (
);

FILL FILL_0__18094_ (
);

FILL FILL432440x93860 (
);

DFFSR _10886_ (
    .CLK(clk_bF$buf83),
    .D(_1191_[11]),
    .Q(\datapath_1.regfile_1.regOut[19] [11]),
    .R(rst_bF$buf81),
    .S(vdd)
);

AND2X2 _10466_ (
    .A(_1042_),
    .B(_1041_),
    .Y(_993_[24])
);

AND2X2 _10046_ (
    .A(_822_),
    .B(_821_),
    .Y(_795_[13])
);

FILL FILL_0__16827_ (
);

FILL FILL_0__16407_ (
);

FILL FILL98800x256880 (
);

FILL FILL_0__11122_ (
);

FILL FILL_0__19299_ (
);

OR2X2 _19164_ (
    .A(_8028_),
    .B(_8062_),
    .Y(_8063_)
);

OR2X2 _8614_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .B(_134__bF$buf0),
    .Y(_88_)
);

FILL FILL345800x24700 (
);

FILL FILL225720x350740 (
);

FILL FILL_1__18619_ (
);

FILL FILL326040x237120 (
);

FILL FILL_0__12747_ (
);

XOR2X1 _12612_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2177_)
);

FILL FILL408880x316160 (
);

AOI22X1 _15084_ (
    .A(_4018_),
    .B(_4013_),
    .C(_4030_),
    .D(_4020_),
    .Y(_4069_)
);

OR2X2 _9819_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_711_)
);

FILL FILL_0__16580_ (
);

FILL FILL_0__16160_ (
);

FILL FILL242440x266760 (
);

FILL FILL_1__14959_ (
);

OR2X2 _13817_ (
    .A(\datapath_1.a [0]),
    .B(_3342__bF$buf3),
    .Y(_3278_)
);

FILL FILL_1__15900_ (
);

AND2X2 _16289_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_5231_)
);

FILL FILL_1__18372_ (
);

FILL FILL288800x83980 (
);

FILL FILL88160x133380 (
);

FILL FILL152760x74100 (
);

OR2X2 _17650_ (
    .A(_6571_),
    .B(_6568_),
    .Y(_6572_)
);

AND2X2 _17230_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_6157_)
);

FILL FILL_0__12080_ (
);

DFFSR _9992_ (
    .CLK(clk_bF$buf44),
    .D(_729_[20]),
    .Q(\datapath_1.regfile_1.regOut[12] [20]),
    .R(rst_bF$buf16),
    .S(vdd)
);

AND2X2 _9572_ (
    .A(_586_),
    .B(_585_),
    .Y(_531_[27])
);

AND2X2 _9152_ (
    .A(_366_),
    .B(_365_),
    .Y(_333_[16])
);

FILL FILL_1__11820_ (
);

FILL FILL_0__10813_ (
);

OR2X2 _18855_ (
    .A(_7750_),
    .B(_7757_),
    .Y(_7758_)
);

FILL FILL_0_BUFX2_insert720 (
);

FILL FILL_0_BUFX2_insert721 (
);

AND2X2 _18435_ (
    .A(_6293__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_7345_)
);

FILL FILL_0_BUFX2_insert722 (
);

OR2X2 _18015_ (
    .A(_6927_),
    .B(_6930_),
    .Y(_6931_)
);

FILL FILL_0_BUFX2_insert723 (
);

OR2X2 _13990_ (
    .A(_3409_),
    .B(_3410_),
    .Y(_3411_)
);

FILL FILL_0__13285_ (
);

FILL FILL_0_BUFX2_insert725 (
);

OR2X2 _13570_ (
    .A(IorD_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [27]),
    .Y(_3068_)
);

OR2X2 _13150_ (
    .A(_2387__bF$buf0),
    .B(_2700_),
    .Y(_2701_)
);

FILL FILL_0_BUFX2_insert727 (
);

FILL FILL_0_BUFX2_insert729 (
);

FILL FILL_0__19511_ (
);

FILL FILL77520x276640 (
);

FILL FILL162640x242060 (
);

FILL FILL136040x207480 (
);

FILL FILL_1__12605_ (
);

FILL FILL223440x212420 (
);

FILL FILL_1__15077_ (
);

FILL FILL117040x365560 (
);

OR2X2 _14775_ (
    .A(\datapath_1.rd2 [6]),
    .B(_3935__bF$buf2),
    .Y(_3883_)
);

DFFSR _14355_ (
    .CLK(clk_bF$buf41),
    .D(_3606_[19]),
    .Q(ALUOut[19]),
    .R(rst_bF$buf63),
    .S(vdd)
);

FILL FILL_0__15851_ (
);

FILL FILL54720x301340 (
);

OR2X2 _10695_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_1155_)
);

FILL FILL_1__17223_ (
);

OR2X2 _10275_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_935_)
);

OR2X2 _16921_ (
    .A(_5852_),
    .B(_5837_),
    .Y(_5853_)
);

FILL FILL_0__16216_ (
);

OR2X2 _16501_ (
    .A(_5439_),
    .B(_5438_),
    .Y(_5440_)
);

FILL FILL_0__11351_ (
);

FILL FILL329840x19760 (
);

AND2X2 _19393_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_8288_)
);

FILL FILL288800x217360 (
);

OR2X2 _8843_ (
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .Y(_265_)
);

BUFX2 _8423_ (
    .A(_1_[31]),
    .Y(memoryAddress[31])
);

FILL FILL_1__18848_ (
);

AND2X2 _17706_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_6627_)
);

FILL FILL_0__12976_ (
);

NOR2X1 _12841_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2406_)
);

FILL FILL_0__12556_ (
);

FILL FILL52440x375440 (
);

FILL FILL_0__12136_ (
);

OR2X2 _12421_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_2048__bF$buf2),
    .Y(_2046_)
);

OR2X2 _12001_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .B(_1850__bF$buf3),
    .Y(_1826_)
);

OR2X2 _9628_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .B(_662__bF$buf2),
    .Y(_604_)
);

DFFSR _9208_ (
    .CLK(clk_bF$buf33),
    .D(_333_[10]),
    .Q(\datapath_1.regfile_1.regOut[6] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

FILL FILL177840x98800 (
);

FILL FILL_1__14768_ (
);

FILL FILL56240x296400 (
);

FILL FILL443080x197600 (
);

AND2X2 _13626_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[5]),
    .Y(_3116_)
);

NAND2X1 _13206_ (
    .A(_2524_),
    .B(_2753_),
    .Y(_2754_)
);

AND2X2 _16098_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_5043_)
);

FILL FILL_0__17594_ (
);

FILL FILL_0__17174_ (
);

FILL FILL126920x256880 (
);

FILL FILL_1__16914_ (
);

OR2X2 _9381_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_479_)
);

FILL FILL_0__10202_ (
);

FILL FILL_0__18799_ (
);

NOR2X1 _18664_ (
    .A(_6310__bF$buf1),
    .B(_7569_),
    .Y(_7570_)
);

FILL FILL_0__18379_ (
);

FILL FILL213560x167960 (
);

AND2X2 _18244_ (
    .A(_6250__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_7157_)
);

FILL FILL_0__19320_ (
);

FILL FILL431680x291460 (
);

FILL FILL281200x24700 (
);

FILL FILL236360x251940 (
);

FILL FILL_1__12414_ (
);

FILL FILL_0__9841_ (
);

FILL FILL_0__11827_ (
);

FILL FILL_0__9001_ (
);

OR2X2 _19449_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8335_)
);

OR2X2 _19029_ (
    .A(_7928_),
    .B(_7929_),
    .Y(_7930_)
);

FILL FILL_0__14299_ (
);

AND2X2 _14584_ (
    .A(_3795_),
    .B(_3794_),
    .Y(_3738_[28])
);

OR2X2 _14164_ (
    .A(MemToReg_bF$buf4),
    .B(ALUOut[7]),
    .Y(_3554_)
);

FILL FILL253840x261820 (
);

FILL FILL_0__15660_ (
);

FILL FILL_0__15240_ (
);

FILL FILL96520x98800 (
);

FILL FILL_1_BUFX2_insert272 (
);

FILL FILL_1_BUFX2_insert274 (
);

FILL FILL_1_BUFX2_insert276 (
);

FILL FILL505400x44460 (
);

AND2X2 _15789_ (
    .A(_4130__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_4739_)
);

OR2X2 _15369_ (
    .A(_4324_),
    .B(_4317_),
    .Y(_4325_)
);

FILL FILL_1__17872_ (
);

OR2X2 _10084_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_860__bF$buf2),
    .Y(_848_)
);

FILL FILL_0__16865_ (
);

AND2X2 _16730_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_5665_)
);

FILL FILL_0__16445_ (
);

FILL FILL_0__16025_ (
);

OR2X2 _16310_ (
    .A(_5251_),
    .B(_5248_),
    .Y(_5252_)
);

FILL FILL471960x251940 (
);

OR2X2 _8652_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_113_)
);

FILL FILL205960x182780 (
);

FILL FILL489440x148200 (
);

FILL FILL_1__18237_ (
);

DFFSR _11289_ (
    .CLK(clk_bF$buf29),
    .D(_1389_[27]),
    .Q(\datapath_1.regfile_1.regOut[22] [27]),
    .R(rst_bF$buf48),
    .S(vdd)
);

AND2X2 _17935_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_6852_)
);

AND2X2 _17515_ (
    .A(_6326__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_6439_)
);

FILL FILL_0__12785_ (
);

FILL FILL_0__12365_ (
);

XNOR2X1 _12650_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2215_)
);

AND2X2 _12230_ (
    .A(_1938_),
    .B(_1937_),
    .Y(_1917_[10])
);

DFFSR _9857_ (
    .CLK(clk_bF$buf3),
    .D(_663_[14]),
    .Q(\datapath_1.regfile_1.regOut[11] [14]),
    .R(rst_bF$buf58),
    .S(vdd)
);

AND2X2 _9437_ (
    .A(_516_),
    .B(_515_),
    .Y(_465_[25])
);

AND2X2 _9017_ (
    .A(_296_),
    .B(_295_),
    .Y(_267_[14])
);

FILL FILL501600x167960 (
);

FILL FILL329840x113620 (
);

FILL FILL35720x39520 (
);

FILL FILL342760x108680 (
);

OR2X2 _13855_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [13]),
    .Y(_3303_)
);

OR2X2 _13435_ (
    .A(_2967_),
    .B(_2376__bF$buf1),
    .Y(_2969_)
);

XOR2X1 _13015_ (
    .A(_2330_),
    .B(_2573_),
    .Y(_2574_)
);

FILL FILL145920x370500 (
);

FILL FILL436240x29640 (
);

FILL FILL_0__14931_ (
);

FILL FILL294120x182780 (
);

FILL FILL23560x276640 (
);

FILL FILL236360x9880 (
);

OR2X2 _9190_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_398__bF$buf4),
    .Y(_392_)
);

FILL FILL_0__15716_ (
);

FILL FILL_1__19195_ (
);

FILL FILL_0__10431_ (
);

FILL FILL_0__10011_ (
);

FILL FILL46360x360620 (
);

OR2X2 _18893_ (
    .A(_7795_),
    .B(_7792_),
    .Y(_7796_)
);

FILL FILL_0__18188_ (
);

AND2X2 _18473_ (
    .A(_6262__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_7382_)
);

AND2X2 _18053_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_6969_)
);

FILL FILL265240x19760 (
);

FILL FILL39520x39520 (
);

FILL FILL363280x266760 (
);

FILL FILL450680x271700 (
);

FILL FILL354920x335920 (
);

FILL FILL_1__12223_ (
);

DFFSR _11921_ (
    .CLK(clk_bF$buf21),
    .D(_1719_[14]),
    .Q(\datapath_1.regfile_1.regOut[27] [14]),
    .R(rst_bF$buf90),
    .S(vdd)
);

FILL FILL_0__11636_ (
);

AND2X2 _11501_ (
    .A(_1572_),
    .B(_1571_),
    .Y(_1521_[25])
);

FILL FILL380760x276640 (
);

OR2X2 _19258_ (
    .A(_8154_),
    .B(_8151_),
    .Y(_8155_)
);

FILL FILL386080x350740 (
);

OR2X2 _14393_ (
    .A(vdd),
    .B(\datapath_1.Data [8]),
    .Y(_3688_)
);

DFFSR _8708_ (
    .CLK(clk_bF$buf55),
    .D(_69_[26]),
    .Q(\datapath_1.regfile_1.regOut[2] [26]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL238640x4940 (
);

FILL FILL_1__13428_ (
);

INVX1 _12706_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .Y(_2271_)
);

FILL FILL142880x93860 (
);

OR2X2 _15598_ (
    .A(_4549_),
    .B(_4550_),
    .Y(_4551_)
);

FILL FILL120080x375440 (
);

AND2X2 _15178_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [0]),
    .Y(_4136_)
);

FILL FILL257640x301340 (
);

FILL FILL_0__16674_ (
);

FILL FILL257640x4940 (
);

FILL FILL329840x340860 (
);

OR2X2 _8881_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_266__bF$buf0),
    .Y(_226_)
);

FILL FILL344280x212420 (
);

OR2X2 _8461_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_68__bF$buf1),
    .Y(_6_)
);

FILL FILL_1__18886_ (
);

OR2X2 _11098_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .B(_1388__bF$buf2),
    .Y(_1364_)
);

FILL FILL_1__13181_ (
);

FILL FILL355680x281580 (
);

FILL FILL_0__17459_ (
);

AND2X2 _17744_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_6664_)
);

FILL FILL_0__17039_ (
);

AND2X2 _17324_ (
    .A(_6249_),
    .B(_6201_),
    .Y(_6250_)
);

FILL FILL_0__18820_ (
);

OR2X2 _9666_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_629_)
);

OR2X2 _9246_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_409_)
);

FILL FILL316160x345800 (
);

FILL FILL192280x123500 (
);

FILL FILL_0__8501_ (
);

OR2X2 _18949_ (
    .A(_7847_),
    .B(_7850_),
    .Y(_7851_)
);

OR2X2 _18529_ (
    .A(_7435_),
    .B(_7436_),
    .Y(_7437_)
);

OR2X2 _18109_ (
    .A(_7022_),
    .B(_7023_),
    .Y(_7024_)
);

FILL FILL_1_BUFX2_insert1031 (
);

FILL FILL_1_BUFX2_insert1033 (
);

FILL FILL_0__13799_ (
);

FILL FILL205200x123500 (
);

FILL FILL_0__13379_ (
);

AND2X2 _13664_ (
    .A(_3087__bF$buf0),
    .B(\datapath_1.ALUResult [10]),
    .Y(_3149_)
);

FILL FILL482600x261820 (
);

FILL FILL_1_BUFX2_insert1035 (
);

INVX1 _13244_ (
    .A(_2789_),
    .Y(\datapath_1.ALUResult [12])
);

FILL FILL227240x49400 (
);

FILL FILL_0__14320_ (
);

FILL FILL216600x192660 (
);

FILL FILL_0__9706_ (
);

DFFSR _14869_ (
    .CLK(clk_bF$buf105),
    .D(_3870_[17]),
    .Q(_2_[17]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL414200x222300 (
);

FILL FILL147440x64220 (
);

AND2X2 _14449_ (
    .A(_3725_),
    .B(_3724_),
    .Y(_3672_[26])
);

OR2X2 _14029_ (
    .A(_3444_),
    .B(_3441_),
    .Y(\datapath_1.alu_1.ALUInB [15])
);

FILL FILL_0__15945_ (
);

FILL FILL_0__15525_ (
);

AND2X2 _15810_ (
    .A(_4151__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_4759_)
);

FILL FILL112480x256880 (
);

OR2X2 _18282_ (
    .A(_7193_),
    .B(_7192_),
    .Y(_7194_)
);

OR2X2 _10789_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .B(_1256__bF$buf4),
    .Y(_1198_)
);

FILL FILL_1__17737_ (
);

FILL FILL_1__17317_ (
);

DFFSR _10369_ (
    .CLK(clk_bF$buf30),
    .D(_927_[10]),
    .Q(\datapath_1.regfile_1.regOut[15] [10]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL135280x340860 (
);

FILL FILL_1__12032_ (
);

FILL FILL_0__11865_ (
);

FILL FILL_0__11445_ (
);

OR2X2 _11730_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_1685_)
);

FILL FILL116280x177840 (
);

FILL FILL53200x128440 (
);

OR2X2 _11310_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_1465_)
);

OR2X2 _19487_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_8360_)
);

AND2X2 _19067_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_7967_)
);

FILL FILL88920x93860 (
);

OR2X2 _8937_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_263_)
);

OR2X2 _8517_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_43_)
);

FILL FILL500080x98800 (
);

FILL FILL65360x93860 (
);

NOR2X1 _12935_ (
    .A(_2163_),
    .B(_2498_),
    .Y(_2499_)
);

FILL FILL_1_BUFX2_insert652 (
);

INVX1 _12515_ (
    .A(_2094_),
    .Y(ALUOp[0])
);

FILL FILL_1_BUFX2_insert654 (
);

FILL FILL_1_BUFX2_insert656 (
);

FILL FILL_1__17490_ (
);

FILL FILL_0__16063_ (
);

FILL FILL133000x311220 (
);

FILL FILL351880x177840 (
);

DFFSR _8690_ (
    .CLK(clk_bF$buf3),
    .D(_69_[8]),
    .Q(\datapath_1.regfile_1.regOut[2] [8]),
    .R(rst_bF$buf4),
    .S(vdd)
);

BUFX2 BUFX2_insert320 (
    .A(_464_),
    .Y(_464__bF$buf2)
);

BUFX2 BUFX2_insert321 (
    .A(_464_),
    .Y(_464__bF$buf1)
);

BUFX2 BUFX2_insert322 (
    .A(_464_),
    .Y(_464__bF$buf0)
);

BUFX2 BUFX2_insert323 (
    .A(_2376_),
    .Y(_2376__bF$buf3)
);

BUFX2 BUFX2_insert324 (
    .A(_2376_),
    .Y(_2376__bF$buf2)
);

OR2X2 _17973_ (
    .A(_6889_),
    .B(_6888_),
    .Y(_6890_)
);

FILL FILL_0__17688_ (
);

FILL FILL51680x187720 (
);

FILL FILL_0__17268_ (
);

BUFX2 BUFX2_insert325 (
    .A(_2376_),
    .Y(_2376__bF$buf1)
);

OR2X2 _17553_ (
    .A(_6475_),
    .B(_6474_),
    .Y(_6476_)
);

BUFX2 BUFX2_insert326 (
    .A(_2376_),
    .Y(_2376__bF$buf0)
);

AND2X2 _17133_ (
    .A(_4225__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_6062_)
);

BUFX2 BUFX2_insert327 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf4 )
);

FILL FILL91200x296400 (
);

BUFX2 BUFX2_insert328 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf3 )
);

BUFX2 BUFX2_insert329 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf2 )
);

FILL FILL231040x291460 (
);

FILL FILL108680x192660 (
);

FILL FILL45600x143260 (
);

OR2X2 _9895_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .B(_794__bF$buf0),
    .Y(_742_)
);

DFFSR _9475_ (
    .CLK(clk_bF$buf60),
    .D(_465_[19]),
    .Q(\datapath_1.regfile_1.regOut[8] [19]),
    .R(rst_bF$buf101),
    .S(vdd)
);

OR2X2 _9055_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .B(_332__bF$buf3),
    .Y(_322_)
);

FILL FILL_1__11723_ (
);

FILL FILL258400x9880 (
);

FILL FILL_0__10716_ (
);

AND2X2 _18758_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_7663_)
);

AND2X2 _18338_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_7249_)
);

AND2X2 _13893_ (
    .A(_3328_),
    .B(_3327_),
    .Y(\datapath_1.alu_1.ALUInA [25])
);

FILL FILL_0__13188_ (
);

INVX1 _13473_ (
    .A(RegDst),
    .Y(_3005_)
);

NAND2X1 _13053_ (
    .A(_2267_),
    .B(_2504_),
    .Y(_2610_)
);

FILL FILL414960x217360 (
);

FILL FILL158840x207480 (
);

FILL FILL385320x133380 (
);

FILL FILL235600x172900 (
);

FILL FILL_0__9515_ (
);

FILL FILL437760x301340 (
);

FILL FILL285000x227240 (
);

OR2X2 _14678_ (
    .A(vdd),
    .B(\datapath_1.a [17]),
    .Y(_3838_)
);

OR2X2 _14258_ (
    .A(vdd),
    .B(ALUOut[6]),
    .Y(_3618_)
);

FILL FILL_1__16341_ (
);

FILL FILL106400x163020 (
);

FILL FILL_0__15334_ (
);

AND2X2 _18091_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_7006_)
);

FILL FILL_1__17966_ (
);

AND2X2 _10598_ (
    .A(_1110_),
    .B(_1109_),
    .Y(_1059_[25])
);

AND2X2 _10178_ (
    .A(_890_),
    .B(_889_),
    .Y(_861_[14])
);

FILL FILL_0__16959_ (
);

FILL FILL_0__16539_ (
);

OR2X2 _16824_ (
    .A(_5742_),
    .B(_5757_),
    .Y(_5758_)
);

AND2X2 _16404_ (
    .A(_4135__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_5344_)
);

FILL FILL_0__11254_ (
);

AND2X2 _19296_ (
    .A(_6206__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_8192_)
);

FILL FILL_0__17900_ (
);

OR2X2 _8746_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .B(_200__bF$buf0),
    .Y(_156_)
);

FILL FILL129200x113620 (
);

FILL FILL11400x217360 (
);

FILL FILL_1__13466_ (
);

FILL FILL_1__13046_ (
);

AND2X2 _17609_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_6531_)
);

OR2X2 _12744_ (
    .A(_2308_),
    .B(_2268_),
    .Y(_2309_)
);

DFFSR _12324_ (
    .CLK(clk_bF$buf7),
    .D(_1917_[30]),
    .Q(\datapath_1.regfile_1.regOut[30] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL_0__13820_ (
);

FILL FILL290320x64220 (
);

FILL FILL_0__16292_ (
);

FILL FILL218880x291460 (
);

AND2X2 _13949_ (
    .A(_3350__bF$buf1),
    .B(_2_[4]),
    .Y(_3376_)
);

FILL FILL364040x153140 (
);

OR2X2 _13529_ (
    .A(ALUOut[13]),
    .B(_3079__bF$buf0),
    .Y(_3041_)
);

AND2X2 _13109_ (
    .A(_2662_),
    .B(_2660_),
    .Y(_2663_)
);

FILL FILL465120x74100 (
);

FILL FILL329080x316160 (
);

FILL FILL381520x163020 (
);

FILL FILL_0__17497_ (
);

AND2X2 _17782_ (
    .A(_6271__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [6]),
    .Y(_6702_)
);

AND2X2 _17362_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_6288_)
);

FILL FILL346560x326040 (
);

FILL FILL58520x182780 (
);

FILL FILL190760x316160 (
);

AND2X2 _9284_ (
    .A(_434_),
    .B(_433_),
    .Y(_399_[17])
);

FILL FILL_1__11112_ (
);

FILL FILL_1__19289_ (
);

FILL FILL_0__10945_ (
);

FILL FILL_0__10525_ (
);

OR2X2 _10810_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_1256__bF$buf0),
    .Y(_1212_)
);

AND2X2 _18987_ (
    .A(_6247__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_7888_)
);

FILL FILL22800x69160 (
);

OR2X2 _18567_ (
    .A(_7473_),
    .B(_7474_),
    .Y(_7475_)
);

AND2X2 _18147_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_7061_)
);

OR2X2 _13282_ (
    .A(_2431_),
    .B(_2501_),
    .Y(_2825_)
);

FILL FILL239400x59280 (
);

FILL FILL55480x227240 (
);

FILL FILL146680x29640 (
);

FILL FILL_0__19223_ (
);

FILL FILL81320x360620 (
);

FILL FILL62320x197600 (
);

DFFSR _14487_ (
    .CLK(clk_bF$buf2),
    .D(_3672_[22]),
    .Q(\datapath_1.Data [22]),
    .R(rst_bF$buf26),
    .S(vdd)
);

OR2X2 _14067_ (
    .A(_3475_),
    .B(_3476_),
    .Y(_3477_)
);

FILL FILL_1__16990_ (
);

FILL FILL_1__16570_ (
);

FILL FILL_0__15563_ (
);

FILL FILL_0__15143_ (
);

FILL FILL_1__17355_ (
);

FILL FILL116280x247000 (
);

FILL FILL146680x158080 (
);

OR2X2 _16633_ (
    .A(_5538_),
    .B(_5569_),
    .Y(_5570_)
);

AND2X2 _16213_ (
    .A(_4189__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_5156_)
);

FILL FILL_0__11483_ (
);

FILL FILL_0__11063_ (
);

AND2X2 _8975_ (
    .A(_268_),
    .B(_331_),
    .Y(_267_[0])
);

DFFSR _8555_ (
    .CLK(clk_bF$buf111),
    .D(_3_[2]),
    .Q(\datapath_1.regfile_1.regOut[1] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

FILL FILL_1__10803_ (
);

FILL FILL_1__13695_ (
);

OR2X2 _17838_ (
    .A(_6753_),
    .B(_6756_),
    .Y(_6757_)
);

AND2X2 _17418_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_6343_)
);

XOR2X1 _12973_ (
    .A(_2360_),
    .B(_2484_),
    .Y(_2535_)
);

FILL FILL_0__12688_ (
);

FILL FILL_0__12268_ (
);

FILL FILL_1__19501_ (
);

OR2X2 _12553_ (
    .A(_2106_),
    .B(ALUOp[1]),
    .Y(_2141_)
);

OR2X2 _12133_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .B(_1916__bF$buf4),
    .Y(_1894_)
);

FILL FILL300200x44460 (
);

FILL FILL405840x24700 (
);

FILL FILL390640x281580 (
);

OR2X2 _13758_ (
    .A(_3229_),
    .B(_3226_),
    .Y(\datapath_1.mux_pcsrc.dout [23])
);

INVX1 _13338_ (
    .A(_2878_),
    .Y(\datapath_1.ALUResult [7])
);

FILL FILL287280x326040 (
);

FILL FILL_0__14834_ (
);

BUFX2 BUFX2_insert700 (
    .A(_2387_),
    .Y(_2387__bF$buf3)
);

BUFX2 BUFX2_insert701 (
    .A(_2387_),
    .Y(_2387__bF$buf2)
);

BUFX2 BUFX2_insert702 (
    .A(_2387_),
    .Y(_2387__bF$buf1)
);

BUFX2 BUFX2_insert703 (
    .A(_2387_),
    .Y(_2387__bF$buf0)
);

BUFX2 BUFX2_insert704 (
    .A(_4151_),
    .Y(_4151__bF$buf4)
);

AND2X2 _17591_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_6514_)
);

BUFX2 BUFX2_insert705 (
    .A(_4151_),
    .Y(_4151__bF$buf3)
);

BUFX2 BUFX2_insert706 (
    .A(_4151_),
    .Y(_4151__bF$buf2)
);

OR2X2 _17171_ (
    .A(_6097_),
    .B(_6098_),
    .Y(_6099_)
);

BUFX2 BUFX2_insert707 (
    .A(_4151_),
    .Y(_4151__bF$buf1)
);

BUFX2 BUFX2_insert708 (
    .A(_4151_),
    .Y(_4151__bF$buf0)
);

BUFX2 BUFX2_insert709 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf4 )
);

FILL FILL294120x296400 (
);

FILL FILL130720x4940 (
);

FILL FILL_1__16206_ (
);

DFFSR _9093_ (
    .CLK(clk_bF$buf105),
    .D(_267_[24]),
    .Q(\datapath_1.regfile_1.regOut[5] [24]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL504640x153140 (
);

FILL FILL348840x83980 (
);

FILL FILL248520x143260 (
);

FILL FILL278160x59280 (
);

OR2X2 _15904_ (
    .A(_4851_),
    .B(_4848_),
    .Y(_4852_)
);

FILL FILL_0__10334_ (
);

FILL FILL31160x143260 (
);

AND2X2 _18796_ (
    .A(_6312__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_7700_)
);

OR2X2 _18376_ (
    .A(_7286_),
    .B(_7285_),
    .Y(_7287_)
);

FILL FILL22800x212420 (
);

AOI21X1 _13091_ (
    .A(_2643_),
    .B(_2645_),
    .C(_2642_),
    .Y(_2646_)
);

FILL FILL231040x29640 (
);

FILL FILL429400x39520 (
);

FILL FILL_0__19452_ (
);

FILL FILL_0__9553_ (
);

FILL FILL_0__11959_ (
);

OR2X2 _11824_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .B(_1784__bF$buf0),
    .Y(_1728_)
);

FILL FILL_0__9133_ (
);

DFFSR _11404_ (
    .CLK(clk_bF$buf63),
    .D(_1455_[13]),
    .Q(\datapath_1.regfile_1.regOut[23] [13]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL_0__11119_ (
);

AND2X2 _14296_ (
    .A(_3643_),
    .B(_3642_),
    .Y(_3606_[18])
);

FILL FILL_0__15792_ (
);

FILL FILL20520x286520 (
);

AND2X2 _12609_ (
    .A(_2173_),
    .B(_2169_),
    .Y(_2174_)
);

FILL FILL457520x0 (
);

FILL FILL_0__16577_ (
);

AND2X2 _16862_ (
    .A(_4167__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_5795_)
);

AND2X2 _16442_ (
    .A(_5381_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [18])
);

FILL FILL_0__16157_ (
);

OR2X2 _16022_ (
    .A(_4966_),
    .B(_4967_),
    .Y(_4968_)
);

FILL FILL178600x44460 (
);

OR2X2 _8784_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_181_)
);

AND2X2 _17647_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_6569_)
);

FILL FILL214320x217360 (
);

AND2X2 _17227_ (
    .A(_4146__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_6154_)
);

FILL FILL301720x222300 (
);

NAND2X1 _12782_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(_2346_),
    .Y(_2347_)
);

FILL FILL_0__12497_ (
);

AND2X2 _12362_ (
    .A(_2006_),
    .B(_2005_),
    .Y(_1983_[11])
);

FILL FILL392160x251940 (
);

FILL FILL_0__18723_ (
);

FILL FILL_0__18303_ (
);

DFFSR _9989_ (
    .CLK(clk_bF$buf109),
    .D(_729_[17]),
    .Q(\datapath_1.regfile_1.regOut[12] [17]),
    .R(rst_bF$buf84),
    .S(vdd)
);

AND2X2 _9569_ (
    .A(_584_),
    .B(_583_),
    .Y(_531_[26])
);

AND2X2 _9149_ (
    .A(_364_),
    .B(_363_),
    .Y(_333_[15])
);

FILL FILL231800x227240 (
);

FILL FILL126160x182780 (
);

FILL FILL_0__8404_ (
);

FILL FILL_0_BUFX2_insert690 (
);

FILL FILL_0_BUFX2_insert692 (
);

FILL FILL_0_BUFX2_insert694 (
);

OR2X2 _13987_ (
    .A(_3408_),
    .B(_3405_),
    .Y(\datapath_1.alu_1.ALUInB [9])
);

FILL FILL_0_BUFX2_insert695 (
);

OR2X2 _13567_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [26]),
    .Y(_3066_)
);

OR2X2 _13147_ (
    .A(_2283_),
    .B(_2449_),
    .Y(_2698_)
);

FILL FILL_0_BUFX2_insert696 (
);

FILL FILL_0_BUFX2_insert697 (
);

FILL FILL_0_BUFX2_insert698 (
);

FILL FILL_0_BUFX2_insert699 (
);

FILL FILL_0__14643_ (
);

FILL FILL_1__16855_ (
);

FILL FILL_1__16435_ (
);

FILL FILL_0__15428_ (
);

AND2X2 _15713_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_4664_)
);

FILL FILL_0__10563_ (
);

FILL FILL_0__10143_ (
);

FILL FILL44080x182780 (
);

OR2X2 _18185_ (
    .A(_7098_),
    .B(_7095_),
    .Y(_7099_)
);

FILL FILL278920x192660 (
);

FILL FILL206720x232180 (
);

FILL FILL_0__19261_ (
);

OR2X2 _16918_ (
    .A(_5848_),
    .B(_5849_),
    .Y(_5850_)
);

FILL FILL106400x326040 (
);

FILL FILL_0__11768_ (
);

FILL FILL_0__9362_ (
);

AND2X2 _11633_ (
    .A(_1640_),
    .B(_1639_),
    .Y(_1587_[26])
);

AND2X2 _11213_ (
    .A(_1420_),
    .B(_1419_),
    .Y(_1389_[15])
);

FILL FILL284240x360620 (
);

FILL FILL275880x237120 (
);

FILL FILL341240x24700 (
);

FILL FILL265240x197600 (
);

FILL FILL_0__15181_ (
);

NAND2X1 _12838_ (
    .A(_2196_),
    .B(_2402_),
    .Y(_2403_)
);

OR2X2 _12418_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .B(_2048__bF$buf4),
    .Y(_2044_)
);

FILL FILL210520x247000 (
);

FILL FILL_1__14921_ (
);

FILL FILL_0__13914_ (
);

FILL FILL193800x14820 (
);

FILL FILL_0__16386_ (
);

OR2X2 _16671_ (
    .A(_5605_),
    .B(_5606_),
    .Y(_5607_)
);

AND2X2 _16251_ (
    .A(_4187__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_5193_)
);

FILL FILL_1__9523_ (
);

FILL FILL491720x83980 (
);

OR2X2 _8593_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .B(_134__bF$buf2),
    .Y(_74_)
);

FILL FILL328320x237120 (
);

FILL FILL_1__18178_ (
);

OR2X2 _17876_ (
    .A(_6793_),
    .B(_6792_),
    .Y(_6794_)
);

OR2X2 _17456_ (
    .A(_6373_),
    .B(_6380_),
    .Y(_6381_)
);

OR2X2 _17036_ (
    .A(_5964_),
    .B(_5965_),
    .Y(_5966_)
);

NAND3X1 _12591_ (
    .A(_2154_),
    .B(ALUControl[1]),
    .C(_2155_),
    .Y(_2156_)
);

DFFSR _12171_ (
    .CLK(clk_bF$buf14),
    .D(_1851_[6]),
    .Q(\datapath_1.regfile_1.regOut[29] [6]),
    .R(rst_bF$buf8),
    .S(vdd)
);

FILL FILL_0__18952_ (
);

OR2X2 _9798_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_697_)
);

FILL FILL244720x266760 (
);

OR2X2 _9378_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_477_)
);

FILL FILL197600x14820 (
);

FILL FILL_0__8633_ (
);

DFFSR _10904_ (
    .CLK(clk_bF$buf6),
    .D(_1191_[29]),
    .Q(\datapath_1.regfile_1.regOut[19] [29]),
    .R(rst_bF$buf31),
    .S(vdd)
);

FILL FILL176320x148200 (
);

OR2X2 _13796_ (
    .A(_3260_),
    .B(_3261_),
    .Y(_3262_)
);

AND2X2 _13376_ (
    .A(_2911_),
    .B(_2913_),
    .Y(_2914_)
);

FILL FILL162640x172900 (
);

FILL FILL_0__19317_ (
);

FILL FILL_0__14452_ (
);

FILL FILL_0__14032_ (
);

FILL FILL_0__9838_ (
);

FILL FILL_0__9418_ (
);

FILL FILL449160x167960 (
);

FILL FILL174800x88920 (
);

AND2X2 _15942_ (
    .A(_4130__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_4889_)
);

FILL FILL_0__15657_ (
);

AND2X2 _15522_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_4476_)
);

AOI21X1 _15102_ (
    .A(_4005_),
    .B(_4017_),
    .C(_4065__bF$buf2),
    .Y(_4084_)
);

FILL FILL485640x340860 (
);

FILL FILL79800x276640 (
);

FILL FILL_0__19070_ (
);

FILL FILL_1__12164_ (
);

FILL FILL119320x365560 (
);

OR2X2 _16727_ (
    .A(_5658_),
    .B(_5661_),
    .Y(_5662_)
);

AND2X2 _16307_ (
    .A(_4181__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_5249_)
);

FILL FILL251560x153140 (
);

FILL FILL_0__11997_ (
);

FILL FILL_0__11577_ (
);

OR2X2 _11862_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_1753_)
);

OR2X2 _11442_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_1533_)
);

DFFSR _11022_ (
    .CLK(clk_bF$buf37),
    .D(_1257_[18]),
    .Q(\datapath_1.regfile_1.regOut[20] [18]),
    .R(rst_bF$buf87),
    .S(vdd)
);

AND2X2 _19199_ (
    .A(_6255__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_8097_)
);

FILL FILL_0__17803_ (
);

OR2X2 _8649_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_111_)
);

FILL FILL380760x98800 (
);

FILL FILL223440x286520 (
);

XNOR2X1 _12647_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2212_)
);

AND2X2 _12227_ (
    .A(_1936_),
    .B(_1935_),
    .Y(_1917_[9])
);

FILL FILL4560x242060 (
);

FILL FILL_1__14310_ (
);

FILL FILL_0__13303_ (
);

FILL FILL443080x108680 (
);

FILL FILL_0_BUFX2_insert1040 (
);

FILL FILL240920x296400 (
);

FILL FILL57000x98800 (
);

FILL FILL_0_BUFX2_insert1041 (
);

FILL FILL_0_BUFX2_insert1042 (
);

OR2X2 _16480_ (
    .A(_5418_),
    .B(_5415_),
    .Y(_5419_)
);

AND2X2 _16060_ (
    .A(_4239__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_5005_)
);

FILL FILL_0_BUFX2_insert1044 (
);

FILL FILL_0_BUFX2_insert1046 (
);

FILL FILL69160x153140 (
);

FILL FILL_0_BUFX2_insert1048 (
);

FILL FILL_1__15935_ (
);

FILL FILL_1__10650_ (
);

FILL FILL_0__14928_ (
);

FILL FILL_0__14508_ (
);

FILL FILL54720x375440 (
);

OR2X2 _17685_ (
    .A(_6605_),
    .B(_6601_),
    .Y(_6606_)
);

AND2X2 _17265_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_6192_)
);

FILL FILL358720x286520 (
);

FILL FILL291080x340860 (
);

FILL FILL384560x98800 (
);

FILL FILL_0__18341_ (
);

FILL FILL249280x34580 (
);

OR2X2 _9187_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .B(_398__bF$buf0),
    .Y(_390_)
);

FILL FILL_1__11855_ (
);

FILL FILL_0__8442_ (
);

FILL FILL_0__10848_ (
);

OR2X2 _10713_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_1167_)
);

AND2X2 _13185_ (
    .A(_2733_),
    .B(_2728_),
    .Y(_2734_)
);

AND2X2 _19411_ (
    .A(_6262__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_8306_)
);

FILL FILL_0__19126_ (
);

FILL FILL_0__14681_ (
);

FILL FILL_0__14261_ (
);

FILL FILL504640x316160 (
);

FILL FILL_0__9647_ (
);

FILL FILL18240x311220 (
);

DFFSR _11918_ (
    .CLK(clk_bF$buf79),
    .D(_1719_[11]),
    .Q(\datapath_1.regfile_1.regOut[27] [11]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL234840x330980 (
);

FILL FILL_0__15886_ (
);

OR2X2 _15751_ (
    .A(_4699_),
    .B(_4700_),
    .Y(_4701_)
);

FILL FILL_0__15046_ (
);

OR2X2 _15331_ (
    .A(_4286_),
    .B(_4287_),
    .Y(_4288_)
);

FILL FILL_0__10181_ (
);

FILL FILL348080x163020 (
);

FILL FILL_1__8603_ (
);

FILL FILL361000x350740 (
);

FILL FILL351880x0 (
);

FILL FILL207480x64220 (
);

FILL FILL288040x306280 (
);

AND2X2 _16956_ (
    .A(_4203__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_5887_)
);

OR2X2 _16536_ (
    .A(_5466_),
    .B(_5473_),
    .Y(_5474_)
);

AND2X2 _16116_ (
    .A(_4177__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_5061_)
);

FILL FILL138320x345800 (
);

DFFSR _11671_ (
    .CLK(clk_bF$buf82),
    .D(_1587_[22]),
    .Q(\datapath_1.regfile_1.regOut[25] [22]),
    .R(rst_bF$buf94),
    .S(vdd)
);

FILL FILL_0__11386_ (
);

OR2X2 _11251_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .B(_1454__bF$buf0),
    .Y(_1446_)
);

FILL FILL_1__9808_ (
);

OR2X2 _8878_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .B(_266__bF$buf4),
    .Y(_224_)
);

OR2X2 _8458_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_68__bF$buf4),
    .Y(_4_)
);

FILL FILL435480x14820 (
);

NOR2X1 _12876_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2441_)
);

INVX1 _12456_ (
    .A(\aluControl_1.inst [4]),
    .Y(_2050_)
);

DFFSR _12036_ (
    .CLK(clk_bF$buf105),
    .D(_1785_[0]),
    .Q(\datapath_1.regfile_1.regOut[28] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

FILL FILL_0__18817_ (
);

FILL FILL_0__13952_ (
);

FILL FILL_0__13532_ (
);

FILL FILL_0__8918_ (
);

FILL FILL_1__15324_ (
);

FILL FILL227240x326040 (
);

FILL FILL_0__14317_ (
);

DFFSR _14602_ (
    .CLK(clk_bF$buf23),
    .D(_3738_[8]),
    .Q(\datapath_1.PCJump [10]),
    .R(rst_bF$buf22),
    .S(vdd)
);

FILL FILL412680x88920 (
);

AND2X2 _17494_ (
    .A(_6262__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_6418_)
);

OR2X2 _17074_ (
    .A(_6002_),
    .B(_6003_),
    .Y(_6004_)
);

FILL FILL_0__18990_ (
);

FILL FILL_0__18570_ (
);

FILL FILL_0__18150_ (
);

FILL FILL439280x14820 (
);

FILL FILL_1__16949_ (
);

FILL FILL_1__11244_ (
);

AND2X2 _15807_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_4756_)
);

FILL FILL_0__8671_ (
);

OR2X2 _10942_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .B(_1322__bF$buf1),
    .Y(_1280_)
);

FILL FILL_0__10657_ (
);

OR2X2 _10522_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(_1124__bF$buf1),
    .Y(_1060_)
);

DFFSR _10102_ (
    .CLK(clk_bF$buf106),
    .D(_795_[1]),
    .Q(\datapath_1.regfile_1.regOut[13] [1]),
    .R(rst_bF$buf96),
    .S(vdd)
);

AND2X2 _18699_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_7605_)
);

INVX1 _18279_ (
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_7191_)
);

AND2X2 _19220_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_8118_)
);

FILL FILL296400x182780 (
);

FILL FILL_0__14070_ (
);

FILL FILL_0__9036_ (
);

OR2X2 _11727_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_1683_)
);

OR2X2 _11307_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_1463_)
);

AND2X2 _14199_ (
    .A(_3577_),
    .B(_3576_),
    .Y(\datapath_1.mux_wd3.dout [18])
);

FILL FILL_0__12803_ (
);

FILL FILL48640x360620 (
);

AND2X2 _15980_ (
    .A(_4239__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_4927_)
);

FILL FILL_0__15695_ (
);

FILL FILL288040x19760 (
);

FILL FILL_0__15275_ (
);

OR2X2 _15560_ (
    .A(_4512_),
    .B(_4509_),
    .Y(_4513_)
);

AND2X2 _15140_ (
    .A(_4108_),
    .B(_4069_),
    .Y(_4109_)
);

FILL FILL_1__8412_ (
);

FILL FILL365560x266760 (
);

FILL FILL388360x350740 (
);

FILL FILL310840x316160 (
);

OR2X2 _16765_ (
    .A(_5697_),
    .B(_5698_),
    .Y(_5699_)
);

OR2X2 _16345_ (
    .A(_5270_),
    .B(_5285_),
    .Y(_5286_)
);

AND2X2 _11480_ (
    .A(_1558_),
    .B(_1557_),
    .Y(_1521_[18])
);

FILL FILL_0__11195_ (
);

AND2X2 _11060_ (
    .A(_1338_),
    .B(_1337_),
    .Y(_1323_[7])
);

FILL FILL_1__9617_ (
);

FILL FILL_0__17841_ (
);

FILL FILL_0__17421_ (
);

DFFSR _8687_ (
    .CLK(clk_bF$buf68),
    .D(_69_[5]),
    .Q(\datapath_1.regfile_1.regOut[2] [5]),
    .R(rst_bF$buf21),
    .S(vdd)
);

FILL FILL_1__10935_ (
);

FILL FILL306280x118560 (
);

BUFX2 BUFX2_insert290 (
    .A(_4181_),
    .Y(_4181__bF$buf2)
);

BUFX2 BUFX2_insert291 (
    .A(_4181_),
    .Y(_4181__bF$buf1)
);

BUFX2 BUFX2_insert292 (
    .A(_4181_),
    .Y(_4181__bF$buf0)
);

BUFX2 BUFX2_insert293 (
    .A(_200_),
    .Y(_200__bF$buf4)
);

BUFX2 BUFX2_insert294 (
    .A(_200_),
    .Y(_200__bF$buf3)
);

BUFX2 BUFX2_insert295 (
    .A(_200_),
    .Y(_200__bF$buf2)
);

BUFX2 BUFX2_insert296 (
    .A(_200_),
    .Y(_200__bF$buf1)
);

BUFX2 BUFX2_insert297 (
    .A(_200_),
    .Y(_200__bF$buf0)
);

FILL FILL122360x375440 (
);

BUFX2 BUFX2_insert298 (
    .A(_3737_),
    .Y(_3737__bF$buf4)
);

AND2X2 _12685_ (
    .A(_2249_),
    .B(_2245_),
    .Y(_2250_)
);

BUFX2 BUFX2_insert299 (
    .A(_3737_),
    .Y(_3737__bF$buf3)
);

OR2X2 _12265_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .B(_1982__bF$buf2),
    .Y(_1962_)
);

OR2X2 _18911_ (
    .A(_7812_),
    .B(_7811_),
    .Y(_7813_)
);

FILL FILL_0__18206_ (
);

FILL FILL418000x266760 (
);

FILL FILL505400x271700 (
);

FILL FILL_0__8727_ (
);

FILL FILL346560x212420 (
);

FILL FILL_1__15973_ (
);

FILL FILL_1__15553_ (
);

FILL FILL_0__14966_ (
);

OR2X2 _14831_ (
    .A(vdd),
    .B(_2_[25]),
    .Y(_3920_)
);

FILL FILL_0__14126_ (
);

OR2X2 _14411_ (
    .A(vdd),
    .B(\datapath_1.Data [14]),
    .Y(_3700_)
);

FILL FILL_1__11053_ (
);

FILL FILL344280x286520 (
);

OR2X2 _15616_ (
    .A(_4566_),
    .B(_4567_),
    .Y(_4568_)
);

FILL FILL_0__10466_ (
);

DFFSR _10751_ (
    .CLK(clk_bF$buf68),
    .D(_1125_[5]),
    .Q(\datapath_1.regfile_1.regOut[18] [5]),
    .R(rst_bF$buf40),
    .S(vdd)
);

AND2X2 _10331_ (
    .A(_972_),
    .B(_971_),
    .Y(_927_[22])
);

OR2X2 _18088_ (
    .A(_7002_),
    .B(_6999_),
    .Y(_7003_)
);

FILL FILL_0__19164_ (
);

FILL FILL_1__12678_ (
);

FILL FILL_0__9685_ (
);

FILL FILL_0__9265_ (
);

OR2X2 _11956_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .B(_1850__bF$buf2),
    .Y(_1796_)
);

FILL FILL354160x64220 (
);

DFFSR _11536_ (
    .CLK(clk_bF$buf76),
    .D(_1521_[16]),
    .Q(\datapath_1.regfile_1.regOut[24] [16]),
    .R(rst_bF$buf112),
    .S(vdd)
);

OR2X2 _11116_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .B(_1388__bF$buf3),
    .Y(_1376_)
);

FILL FILL192280x197600 (
);

FILL FILL_0__12612_ (
);

FILL FILL410400x375440 (
);

FILL FILL_0__15084_ (
);

FILL FILL341240x182780 (
);

FILL FILL137560x340860 (
);

FILL FILL_1__17296_ (
);

AND2X2 _16994_ (
    .A(_4142__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_5925_)
);

AND2X2 _16574_ (
    .A(_4158__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_5511_)
);

AND2X2 _16154_ (
    .A(_4158__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_5098_)
);

OR2X2 _8496_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_29_)
);

FILL FILL_1__10744_ (
);

FILL FILL241680x261820 (
);

FILL FILL88160x93860 (
);

FILL FILL281200x370500 (
);

FILL FILL395200x118560 (
);

OR2X2 _17779_ (
    .A(_6697_),
    .B(_6698_),
    .Y(_6699_)
);

FILL FILL448400x9880 (
);

AND2X2 _17359_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_6285_)
);

AND2X2 _12494_ (
    .A(_2095_),
    .B(_2096_),
    .Y(ALUOp[1])
);

AND2X2 _12074_ (
    .A(_1854_),
    .B(_1853_),
    .Y(_1851_[1])
);

FILL FILL_0__18855_ (
);

AND2X2 _18720_ (
    .A(_6259__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_7625_)
);

FILL FILL_0__18435_ (
);

FILL FILL376200x276640 (
);

OR2X2 _18300_ (
    .A(_7208_),
    .B(_7211_),
    .Y(_7212_)
);

FILL FILL_0__18015_ (
);

FILL FILL_0__13570_ (
);

FILL FILL_0__13150_ (
);

FILL FILL212800x9880 (
);

FILL FILL298680x281580 (
);

FILL FILL_0__8536_ (
);

OR2X2 _10807_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_1256__bF$buf4),
    .Y(_1210_)
);

FILL FILL399000x360620 (
);

FILL FILL72960x350740 (
);

AND2X2 _13699_ (
    .A(_3087__bF$buf0),
    .B(\datapath_1.ALUResult [15]),
    .Y(_3179_)
);

XOR2X1 _13279_ (
    .A(_2229_),
    .B(_2821_),
    .Y(_2822_)
);

OR2X2 _19505_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [26]),
    .Y(_8372_)
);

FILL FILL289560x256880 (
);

FILL FILL_0__14775_ (
);

OR2X2 _14640_ (
    .A(\datapath_1.rd1 [4]),
    .B(_3869__bF$buf4),
    .Y(_3813_)
);

AND2X2 _14220_ (
    .A(_3591_),
    .B(_3590_),
    .Y(\datapath_1.mux_wd3.dout [25])
);

FILL FILL233320x291460 (
);

FILL FILL212800x34580 (
);

AND2X2 _15845_ (
    .A(_4200__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_4794_)
);

OR2X2 _15425_ (
    .A(_4376_),
    .B(_4379_),
    .Y(_4380_)
);

DFFSR _15005_ (
    .CLK(clk_bF$buf20),
    .D(_3936_[24]),
    .Q(\datapath_1.mux_iord.din0 [24]),
    .R(rst_bF$buf29),
    .S(vdd)
);

FILL FILL110960x286520 (
);

FILL FILL_0__10695_ (
);

OR2X2 _10980_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_1305_)
);

OR2X2 _10560_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_1085_)
);

FILL FILL_0__10275_ (
);

OR2X2 _10140_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_865_)
);

FILL FILL_0__16921_ (
);

FILL FILL317680x113620 (
);

FILL FILL387600x133380 (
);

FILL FILL_0__19393_ (
);

FILL FILL_0__9494_ (
);

FILL FILL_1__18713_ (
);

AND2X2 _11765_ (
    .A(_1708_),
    .B(_1707_),
    .Y(_1653_[27])
);

AND2X2 _11345_ (
    .A(_1488_),
    .B(_1487_),
    .Y(_1455_[16])
);

FILL FILL_0__17706_ (
);

FILL FILL_0__12001_ (
);

FILL FILL121600x158080 (
);

FILL FILL370880x202540 (
);

OR2X2 _9913_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .B(_794__bF$buf2),
    .Y(_754_)
);

FILL FILL332880x197600 (
);

AND2X2 _13911_ (
    .A(_3340_),
    .B(_3339_),
    .Y(\datapath_1.alu_1.ALUInA [31])
);

FILL FILL_0__13626_ (
);

FILL FILL281960x365560 (
);

AND2X2 _16383_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_5323_)
);

FILL FILL_0__16098_ (
);

FILL FILL_1__9655_ (
);

FILL FILL_1__15418_ (
);

FILL FILL_1__10553_ (
);

BUFX2 BUFX2_insert670 (
    .A(_3081_),
    .Y(_3081__bF$buf4)
);

BUFX2 BUFX2_insert671 (
    .A(_3081_),
    .Y(_3081__bF$buf3)
);

BUFX2 BUFX2_insert672 (
    .A(_3081_),
    .Y(_3081__bF$buf2)
);

BUFX2 BUFX2_insert673 (
    .A(_3081_),
    .Y(_3081__bF$buf1)
);

BUFX2 BUFX2_insert674 (
    .A(_3081_),
    .Y(_3081__bF$buf0)
);

AND2X2 _17588_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_6511_)
);

BUFX2 BUFX2_insert675 (
    .A(_992_),
    .Y(_992__bF$buf4)
);

BUFX2 BUFX2_insert676 (
    .A(_992_),
    .Y(_992__bF$buf3)
);

OR2X2 _17168_ (
    .A(_6092_),
    .B(_6095_),
    .Y(_6096_)
);

BUFX2 BUFX2_insert677 (
    .A(_992_),
    .Y(_992__bF$buf2)
);

BUFX2 BUFX2_insert678 (
    .A(_992_),
    .Y(_992__bF$buf1)
);

FILL FILL91200x345800 (
);

BUFX2 BUFX2_insert679 (
    .A(_992_),
    .Y(_992__bF$buf0)
);

FILL FILL_0__18664_ (
);

FILL FILL_0__18244_ (
);

FILL FILL129200x187720 (
);

AND2X2 _10616_ (
    .A(_1122_),
    .B(_1121_),
    .Y(_1059_[31])
);

FILL FILL101840x49400 (
);

NAND2X1 _13088_ (
    .A(ALUControl[1]),
    .B(_2467_),
    .Y(_2643_)
);

FILL FILL266000x247000 (
);

FILL FILL_0__19029_ (
);

AND2X2 _19314_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_8210_)
);

FILL FILL_0__14584_ (
);

FILL FILL348840x326040 (
);

FILL FILL252320x271700 (
);

FILL FILL_1__16376_ (
);

FILL FILL62320x19760 (
);

FILL FILL_0__15369_ (
);

OR2X2 _15654_ (
    .A(_4604_),
    .B(_4605_),
    .Y(_4606_)
);

OR2X2 _15234_ (
    .A(_4185_),
    .B(_4191_),
    .Y(_4192_)
);

FILL FILL_0__10084_ (
);

FILL FILL_1__8506_ (
);

FILL FILL_0__16310_ (
);

FILL FILL47120x187720 (
);

FILL FILL383040x256880 (
);

FILL FILL83600x360620 (
);

FILL FILL470440x261820 (
);

FILL FILL64600x197600 (
);

AND2X2 _16859_ (
    .A(_4158__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_5792_)
);

OR2X2 _16439_ (
    .A(_5378_),
    .B(_5371_),
    .Y(_5379_)
);

OR2X2 _16019_ (
    .A(_4964_),
    .B(_4963_),
    .Y(_4965_)
);

OR2X2 _11994_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_1821_)
);

OR2X2 _11574_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_1601_)
);

DFFSR _11154_ (
    .CLK(clk_bF$buf21),
    .D(_1323_[21]),
    .Q(\datapath_1.regfile_1.regOut[21] [21]),
    .R(rst_bF$buf90),
    .S(vdd)
);

FILL FILL_0__17935_ (
);

FILL FILL_0__17515_ (
);

AND2X2 _17800_ (
    .A(_6719_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd1 [6])
);

FILL FILL_0__12650_ (
);

DFFSR _9722_ (
    .CLK(clk_bF$buf22),
    .D(_597_[8]),
    .Q(\datapath_1.regfile_1.regOut[10] [8]),
    .R(rst_bF$buf7),
    .S(vdd)
);

AND2X2 _9302_ (
    .A(_446_),
    .B(_445_),
    .Y(_399_[23])
);

FILL FILL66120x19760 (
);

INVX1 _12779_ (
    .A(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2344_)
);

AND2X2 _12359_ (
    .A(_2004_),
    .B(_2003_),
    .Y(_1983_[10])
);

FILL FILL118560x247000 (
);

FILL FILL148960x158080 (
);

FILL FILL_1__14442_ (
);

FILL FILL_0__13435_ (
);

AND2X2 _13720_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [18]),
    .Y(_3197_)
);

AOI21X1 _13300_ (
    .A(_2424_),
    .B(_2593_),
    .C(_2841_),
    .Y(_2842_)
);

FILL FILL_0__13015_ (
);

FILL FILL44080x79040 (
);

FILL FILL158080x9880 (
);

OR2X2 _16192_ (
    .A(_5133_),
    .B(_5134_),
    .Y(_5135_)
);

OR2X2 _14925_ (
    .A(\datapath_1.mux_pcsrc.dout [13]),
    .B(_4001__bF$buf2),
    .Y(_3963_)
);

OR2X2 _14505_ (
    .A(memoryOutData[2]),
    .B(_3803__bF$buf2),
    .Y(_3743_)
);

AND2X2 _17397_ (
    .A(_6228_),
    .B(\datapath_1.PCJump_27_bF$buf1 ),
    .Y(_6323_)
);

FILL FILL440800x79040 (
);

FILL FILL428640x24700 (
);

FILL FILL_1__19060_ (
);

FILL FILL_0__18893_ (
);

FILL FILL462080x182780 (
);

FILL FILL344280x83980 (
);

FILL FILL81320x222300 (
);

FILL FILL405080x24700 (
);

FILL FILL_1__11987_ (
);

OR2X2 _10845_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_1235_)
);

OR2X2 _10425_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_1015_)
);

INVX2 _10005_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .Y(_860_)
);

FILL FILL289560x326040 (
);

FILL FILL196080x9880 (
);

DFFSR _19543_ (
    .CLK(clk_bF$buf9),
    .D(_8320_[20]),
    .Q(\datapath_1.regfile_1.regOut[0] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

FILL FILL_0__19258_ (
);

OR2X2 _19123_ (
    .A(_8021_),
    .B(_8020_),
    .Y(_8022_)
);

FILL FILL_0__14393_ (
);

FILL FILL256880x187720 (
);

FILL FILL_0__9779_ (
);

FILL FILL_0__9359_ (
);

FILL FILL277400x29640 (
);

FILL FILL461320x29640 (
);

FILL FILL167960x49400 (
);

FILL FILL_0__15598_ (
);

AND2X2 _15883_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_4831_)
);

OR2X2 _15463_ (
    .A(_4414_),
    .B(_4417_),
    .Y(_4418_)
);

NAND3X1 _15043_ (
    .A(_4031_),
    .B(_4017_),
    .C(_4030_),
    .Y(_4032_)
);

FILL FILL186200x316160 (
);

OR2X2 _16668_ (
    .A(_5603_),
    .B(_5602_),
    .Y(_5604_)
);

OR2X2 _16248_ (
    .A(_5190_),
    .B(_5175_),
    .Y(_5191_)
);

FILL FILL_0__11098_ (
);

OR2X2 _11383_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .B(_1520__bF$buf0),
    .Y(_1514_)
);

FILL FILL_0__17324_ (
);

FILL FILL_1__10838_ (
);

FILL FILL326800x197600 (
);

OR2X2 _9951_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_779_)
);

OR2X2 _9531_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_559_)
);

OR2X2 _9111_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_339_)
);

INVX1 _12588_ (
    .A(ALUControl[2]),
    .Y(_2153_)
);

DFFSR _12168_ (
    .CLK(clk_bF$buf10),
    .D(_1851_[3]),
    .Q(\datapath_1.regfile_1.regOut[29] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

AND2X2 _18814_ (
    .A(_6302__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_7718_)
);

FILL FILL_0__18529_ (
);

FILL FILL_0__18109_ (
);

FILL FILL_0_BUFX2_insert311 (
);

FILL FILL_0_BUFX2_insert313 (
);

FILL FILL_0__13664_ (
);

FILL FILL_0_BUFX2_insert315 (
);

FILL FILL_0__13244_ (
);

FILL FILL_0_BUFX2_insert316 (
);

FILL FILL_0_BUFX2_insert317 (
);

FILL FILL_0_BUFX2_insert318 (
);

FILL FILL_0_BUFX2_insert319 (
);

FILL FILL385320x44460 (
);

FILL FILL371640x167960 (
);

FILL FILL9120x9880 (
);

DFFSR _14734_ (
    .CLK(clk_bF$buf38),
    .D(_3804_[11]),
    .Q(\datapath_1.a [11]),
    .R(rst_bF$buf15),
    .S(vdd)
);

AND2X2 _14314_ (
    .A(_3655_),
    .B(_3654_),
    .Y(_3606_[24])
);

FILL FILL_0__15810_ (
);

FILL FILL128440x182780 (
);

FILL FILL_0__18282_ (
);

FILL FILL63080x49400 (
);

AND2X2 _15939_ (
    .A(_4234__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_4886_)
);

OR2X2 _15519_ (
    .A(_4471_),
    .B(_4472_),
    .Y(_4473_)
);

FILL FILL_0__10789_ (
);

OR2X2 _10654_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_1190__bF$buf3),
    .Y(_1128_)
);

FILL FILL_1__17602_ (
);

DFFSR _10234_ (
    .CLK(clk_bF$buf24),
    .D(_861_[4]),
    .Q(\datapath_1.regfile_1.regOut[14] [4]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_0__11730_ (
);

FILL FILL307040x370500 (
);

FILL FILL_0__19487_ (
);

AND2X2 _19352_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_8248_)
);

OR2X2 _8802_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_193_)
);

FILL FILL151240x360620 (
);

FILL FILL142880x237120 (
);

FILL FILL_0__9168_ (
);

OR2X2 _11859_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_1751_)
);

FILL FILL352640x113620 (
);

OR2X2 _11439_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_1531_)
);

DFFSR _11019_ (
    .CLK(clk_bF$buf111),
    .D(_1257_[15]),
    .Q(\datapath_1.regfile_1.regOut[20] [15]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL136040x74100 (
);

FILL FILL_1__13942_ (
);

FILL FILL269800x123500 (
);

INVX1 _12800_ (
    .A(_2356_),
    .Y(_2365_)
);

FILL FILL_0__12515_ (
);

OR2X2 _15692_ (
    .A(_4642_),
    .B(_4641_),
    .Y(_4643_)
);

AND2X2 _15272_ (
    .A(_4216_),
    .B(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_4230_)
);

FILL FILL487160x153140 (
);

FILL FILL117800x59280 (
);

FILL FILL286520x360620 (
);

OR2X2 _16897_ (
    .A(_5825_),
    .B(_5828_),
    .Y(_5829_)
);

AND2X2 _16477_ (
    .A(_4187__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_5416_)
);

OR2X2 _16057_ (
    .A(_4971_),
    .B(_5002_),
    .Y(_5003_)
);

AND2X2 _11192_ (
    .A(_1406_),
    .B(_1405_),
    .Y(_1389_[8])
);

FILL FILL_1__9749_ (
);

FILL FILL_0__17973_ (
);

FILL FILL_0__17553_ (
);

FILL FILL_0__17133_ (
);

BUFX2 _8399_ (
    .A(_1_[7]),
    .Y(memoryAddress[7])
);

FILL FILL277400x335920 (
);

OR2X2 _9760_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .B(_728__bF$buf3),
    .Y(_672_)
);

DFFSR _9340_ (
    .CLK(clk_bF$buf103),
    .D(_399_[13]),
    .Q(\datapath_1.regfile_1.regOut[7] [13]),
    .R(rst_bF$buf32),
    .S(vdd)
);

FILL FILL12920x44460 (
);

OR2X2 _12397_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .B(_2048__bF$buf2),
    .Y(_2030_)
);

FILL FILL_0__18758_ (
);

AND2X2 _18623_ (
    .A(_6236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_7530_)
);

OR2X2 _18203_ (
    .A(_7115_),
    .B(_7114_),
    .Y(_7116_)
);

FILL FILL_0__13893_ (
);

FILL FILL_0__13473_ (
);

FILL FILL_0__13053_ (
);

FILL FILL193040x14820 (
);

FILL FILL_0__8859_ (
);

FILL FILL_0__8439_ (
);

FILL FILL_0__9800_ (
);

FILL FILL116280x69160 (
);

FILL FILL500080x138320 (
);

AND2X2 _19408_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_8303_)
);

OR2X2 _14963_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [26]),
    .Y(_3988_)
);

OR2X2 _14543_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3768_)
);

OR2X2 _14123_ (
    .A(_3523_),
    .B(_3524_),
    .Y(_3525_)
);

FILL FILL12160x256880 (
);

FILL FILL16720x271700 (
);

FILL FILL368600x98800 (
);

OR2X2 _15748_ (
    .A(_4697_),
    .B(_4696_),
    .Y(_4698_)
);

OR2X2 _15328_ (
    .A(_4281_),
    .B(_4284_),
    .Y(_4285_)
);

FILL FILL284240x222300 (
);

DFFSR _10883_ (
    .CLK(clk_bF$buf84),
    .D(_1191_[8]),
    .Q(\datapath_1.regfile_1.regOut[19] [8]),
    .R(rst_bF$buf11),
    .S(vdd)
);

FILL FILL_0__10598_ (
);

FILL FILL_1__17831_ (
);

AND2X2 _10463_ (
    .A(_1040_),
    .B(_1039_),
    .Y(_993_[23])
);

AND2X2 _10043_ (
    .A(_820_),
    .B(_819_),
    .Y(_795_[12])
);

FILL FILL198360x74100 (
);

FILL FILL_0__16824_ (
);

FILL FILL_0__16404_ (
);

FILL FILL129960x335920 (
);

FILL FILL_0__19296_ (
);

OR2X2 _19161_ (
    .A(_8059_),
    .B(_8052_),
    .Y(_8060_)
);

OR2X2 _8611_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .B(_134__bF$buf1),
    .Y(_86_)
);

FILL FILL_0__9397_ (
);

DFFSR _11668_ (
    .CLK(clk_bF$buf81),
    .D(_1587_[19]),
    .Q(\datapath_1.regfile_1.regOut[25] [19]),
    .R(rst_bF$buf19),
    .S(vdd)
);

OR2X2 _11248_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .B(_1454__bF$buf1),
    .Y(_1444_)
);

FILL FILL_0__17609_ (
);

FILL FILL_0__12744_ (
);

FILL FILL310840x202540 (
);

AND2X2 _15081_ (
    .A(_4048_),
    .B(_4066_),
    .Y(_4067_)
);

FILL FILL96520x148200 (
);

OR2X2 _9816_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_709_)
);

FILL FILL_1__14116_ (
);

FILL FILL422560x158080 (
);

FILL FILL_0__13949_ (
);

OR2X2 _13814_ (
    .A(_3277_),
    .B(_3274_),
    .Y(\datapath_1.mux_pcsrc.dout [31])
);

FILL FILL47880x335920 (
);

FILL FILL253840x153140 (
);

FILL FILL_0__13109_ (
);

AND2X2 _16286_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_5228_)
);

FILL FILL218880x316160 (
);

FILL FILL_1__9558_ (
);

FILL FILL_0__17782_ (
);

FILL FILL_0__17362_ (
);

FILL FILL51680x44460 (
);

FILL FILL411920x54340 (
);

FILL FILL225720x286520 (
);

FILL FILL_1__19154_ (
);

FILL FILL204440x54340 (
);

FILL FILL_0__10810_ (
);

AND2X2 _18852_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_7755_)
);

FILL FILL_0__18147_ (
);

AND2X2 _18432_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_7342_)
);

AND2X2 _18012_ (
    .A(_6247__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_6928_)
);

FILL FILL276640x103740 (
);

FILL FILL133000x133380 (
);

FILL FILL449920x123500 (
);

FILL FILL_0__8668_ (
);

OR2X2 _10939_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .B(_1322__bF$buf4),
    .Y(_1278_)
);

DFFSR _10519_ (
    .CLK(clk_bF$buf56),
    .D(_993_[31]),
    .Q(\datapath_1.regfile_1.regOut[16] [31]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL_1__15494_ (
);

FILL FILL479560x34580 (
);

OR2X2 _19217_ (
    .A(_8114_),
    .B(_8113_),
    .Y(_8115_)
);

OR2X2 _14772_ (
    .A(\datapath_1.rd2 [5]),
    .B(_3935__bF$buf0),
    .Y(_3881_)
);

FILL FILL_0__14067_ (
);

DFFSR _14352_ (
    .CLK(clk_bF$buf12),
    .D(_3606_[16]),
    .Q(ALUOut[16]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL31920x14820 (
);

FILL FILL_1__13807_ (
);

AND2X2 _15977_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_4924_)
);

AND2X2 _15557_ (
    .A(_4146__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_4510_)
);

NOR2X1 _15137_ (
    .A(_4022_),
    .B(_4042_),
    .Y(\datapath_1.regfile_1.regEn [20])
);

OR2X2 _10692_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_1153_)
);

OR2X2 _10272_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_933_)
);

FILL FILL_0__16633_ (
);

OR2X2 _19390_ (
    .A(_8284_),
    .B(_8270_),
    .Y(_8285_)
);

DFFSR _8840_ (
    .CLK(clk_bF$buf88),
    .D(_135_[29]),
    .Q(\datapath_1.regfile_1.regOut[3] [29]),
    .R(rst_bF$buf37),
    .S(vdd)
);

BUFX2 _8420_ (
    .A(_1_[28]),
    .Y(memoryAddress[28])
);

FILL FILL420280x207480 (
);

AND2X2 _11897_ (
    .A(_1776_),
    .B(_1775_),
    .Y(_1719_[28])
);

AND2X2 _11477_ (
    .A(_1556_),
    .B(_1555_),
    .Y(_1521_[17])
);

AND2X2 _11057_ (
    .A(_1336_),
    .B(_1335_),
    .Y(_1323_[6])
);

FILL FILL_1__18005_ (
);

FILL FILL_1__13560_ (
);

FILL FILL_0__17838_ (
);

AND2X2 _17703_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_6624_)
);

FILL FILL_0__12133_ (
);

OR2X2 _9625_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .B(_662__bF$buf2),
    .Y(_602_)
);

DFFSR _9205_ (
    .CLK(clk_bF$buf112),
    .D(_333_[7]),
    .Q(\datapath_1.regfile_1.regOut[6] [7]),
    .R(rst_bF$buf3),
    .S(vdd)
);

OR2X2 _18908_ (
    .A(_7809_),
    .B(_7808_),
    .Y(_7810_)
);

FILL FILL386080x242060 (
);

FILL FILL_0__13758_ (
);

AND2X2 _13623_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3114_)
);

FILL FILL_0__13338_ (
);

AND2X2 _13203_ (
    .A(_2751_),
    .B(_2736_),
    .Y(_2752_)
);

OR2X2 _16095_ (
    .A(_5038_),
    .B(_5039_),
    .Y(_5040_)
);

FILL FILL_1__9367_ (
);

FILL FILL272080x360620 (
);

FILL FILL57760x24700 (
);

FILL FILL_1__10685_ (
);

FILL FILL386080x108680 (
);

OR2X2 _14828_ (
    .A(vdd),
    .B(_2_[24]),
    .Y(_3918_)
);

OR2X2 _14408_ (
    .A(vdd),
    .B(\datapath_1.Data [13]),
    .Y(_3698_)
);

FILL FILL253080x197600 (
);

FILL FILL_0__15904_ (
);

FILL FILL503120x163020 (
);

FILL FILL_0__18796_ (
);

AND2X2 _18661_ (
    .A(_6293__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_7567_)
);

FILL FILL_0__18376_ (
);

AND2X2 _18241_ (
    .A(_6293__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_7154_)
);

FILL FILL_0__13091_ (
);

FILL FILL_0__8477_ (
);

DFFSR _10748_ (
    .CLK(clk_bF$buf18),
    .D(_1125_[2]),
    .Q(\datapath_1.regfile_1.regOut[18] [2]),
    .R(rst_bF$buf107),
    .S(vdd)
);

AND2X2 _10328_ (
    .A(_970_),
    .B(_969_),
    .Y(_927_[21])
);

FILL FILL_0__11824_ (
);

OR2X2 _19446_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8333_)
);

OR2X2 _19026_ (
    .A(_7925_),
    .B(_7926_),
    .Y(_7927_)
);

AND2X2 _14581_ (
    .A(_3793_),
    .B(_3792_),
    .Y(_3738_[27])
);

OR2X2 _14161_ (
    .A(MemToReg_bF$buf0),
    .B(ALUOut[6]),
    .Y(_3552_)
);

FILL FILL388360x197600 (
);

FILL FILL177840x143260 (
);

FILL FILL342000x370500 (
);

FILL FILL_0__12609_ (
);

FILL FILL_1_BUFX2_insert247 (
);

FILL FILL190760x0 (
);

FILL FILL_1_BUFX2_insert249 (
);

AND2X2 _15786_ (
    .A(_4172__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_4736_)
);

AND2X2 _15366_ (
    .A(_4203__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_4322_)
);

OR2X2 _10081_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .B(_860__bF$buf2),
    .Y(_846_)
);

FILL FILL_1__8638_ (
);

FILL FILL269040x326040 (
);

FILL FILL418000x49400 (
);

FILL FILL_0__16442_ (
);

FILL FILL_0__16022_ (
);

FILL FILL395960x133380 (
);

FILL FILL456760x103740 (
);

FILL FILL_1__18654_ (
);

DFFSR _11286_ (
    .CLK(clk_bF$buf8),
    .D(_1389_[24]),
    .Q(\datapath_1.regfile_1.regOut[22] [24]),
    .R(rst_bF$buf6),
    .S(vdd)
);

FILL FILL437760x261820 (
);

AND2X2 _17932_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_6849_)
);

FILL FILL_0__17647_ (
);

FILL FILL_0__17227_ (
);

OR2X2 _17512_ (
    .A(_6435_),
    .B(_6434_),
    .Y(_6436_)
);

FILL FILL496280x79040 (
);

FILL FILL_0__12782_ (
);

FILL FILL281960x251940 (
);

DFFSR _9854_ (
    .CLK(clk_bF$buf71),
    .D(_663_[11]),
    .Q(\datapath_1.regfile_1.regOut[11] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

AND2X2 _9434_ (
    .A(_514_),
    .B(_513_),
    .Y(_465_[24])
);

AND2X2 _9014_ (
    .A(_294_),
    .B(_293_),
    .Y(_267_[13])
);

FILL FILL458280x0 (
);

FILL FILL_1__19019_ (
);

OR2X2 _18717_ (
    .A(_7620_),
    .B(_7621_),
    .Y(_7622_)
);

FILL FILL454480x177840 (
);

FILL FILL_0__13987_ (
);

FILL FILL281960x24700 (
);

OR2X2 _13852_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [12]),
    .Y(_3301_)
);

FILL FILL_0__13567_ (
);

OR2X2 _13432_ (
    .A(_2964_),
    .B(_2965_),
    .Y(_2966_)
);

INVX1 _13012_ (
    .A(_2571_),
    .Y(\datapath_1.ALUResult [26])
);

FILL FILL213560x212420 (
);

FILL FILL_1__15359_ (
);

FILL FILL5320x93860 (
);

FILL FILL_1__10074_ (
);

OR2X2 _14637_ (
    .A(\datapath_1.rd1 [3]),
    .B(_3869__bF$buf1),
    .Y(_3811_)
);

FILL FILL124640x375440 (
);

AND2X2 _14217_ (
    .A(_3589_),
    .B(_3588_),
    .Y(\datapath_1.mux_wd3.dout [24])
);

FILL FILL_1__16720_ (
);

FILL FILL_1__16300_ (
);

FILL FILL269040x49400 (
);

AND2X2 _18890_ (
    .A(_6229__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_7793_)
);

OR2X2 _18470_ (
    .A(_7376_),
    .B(_7378_),
    .Y(_7379_)
);

AND2X2 _18050_ (
    .A(_6323__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_6966_)
);

FILL FILL348840x212420 (
);

FILL FILL_1__11699_ (
);

FILL FILL70680x242060 (
);

FILL FILL338200x172900 (
);

OR2X2 _10977_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_1303_)
);

OR2X2 _10557_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_1083_)
);

OR2X2 _10137_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_863_)
);

FILL FILL351120x167960 (
);

FILL FILL_0__16918_ (
);

FILL FILL374680x153140 (
);

FILL FILL342760x365560 (
);

FILL FILL_0__11213_ (
);

AND2X2 _19255_ (
    .A(_6247__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_8152_)
);

OR2X2 _14390_ (
    .A(vdd),
    .B(\datapath_1.Data [7]),
    .Y(_3686_)
);

DFFSR _8705_ (
    .CLK(clk_bF$buf45),
    .D(_69_[23]),
    .Q(\datapath_1.regfile_1.regOut[2] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL42560x375440 (
);

FILL FILL173280x266760 (
);

FILL FILL346560x286520 (
);

FILL FILL_0__12838_ (
);

OR2X2 _12703_ (
    .A(_2267_),
    .B(_2264_),
    .Y(_2268_)
);

FILL FILL_0__12418_ (
);

FILL FILL127680x34580 (
);

FILL FILL190760x276640 (
);

OR2X2 _15595_ (
    .A(_4546_),
    .B(_4547_),
    .Y(_4548_)
);

AND2X2 _15175_ (
    .A(_4132_),
    .B(\datapath_1.PCJump [19]),
    .Y(_4133_)
);

FILL FILL_1__8447_ (
);

FILL FILL414200x207480 (
);

FILL FILL_0__16251_ (
);

FILL FILL501600x212420 (
);

AND2X2 _13908_ (
    .A(_3338_),
    .B(_3337_),
    .Y(\datapath_1.alu_1.ALUInA [30])
);

OR2X2 _11095_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_1388__bF$buf4),
    .Y(_1362_)
);

FILL FILL_1__18043_ (
);

FILL FILL4560x335920 (
);

FILL FILL_0__17876_ (
);

OR2X2 _17741_ (
    .A(_6660_),
    .B(_6659_),
    .Y(_6661_)
);

AND2X2 _17321_ (
    .A(_6246_),
    .B(_6201_),
    .Y(_6247_)
);

FILL FILL_0__12591_ (
);

OR2X2 _9663_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_627_)
);

OR2X2 _9243_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_407_)
);

FILL FILL139840x340860 (
);

AND2X2 _18946_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_7848_)
);

INVX1 _18526_ (
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_7434_)
);

FILL FILL340480x227240 (
);

OR2X2 _18106_ (
    .A(_7013_),
    .B(_7020_),
    .Y(_7021_)
);

AND2X2 _13661_ (
    .A(_3081__bF$buf1),
    .B(ALUOut[10]),
    .Y(_3146_)
);

OR2X2 _13241_ (
    .A(_2387__bF$buf3),
    .B(_2786_),
    .Y(_2787_)
);

FILL FILL_1_BUFX2_insert1007 (
);

FILL FILL266000x360620 (
);

FILL FILL_1_BUFX2_insert1009 (
);

FILL FILL34960x256880 (
);

DFFSR _14866_ (
    .CLK(clk_bF$buf58),
    .D(_3870_[14]),
    .Q(_2_[14]),
    .R(rst_bF$buf15),
    .S(vdd)
);

AND2X2 _14446_ (
    .A(_3723_),
    .B(_3722_),
    .Y(_3672_[25])
);

AND2X2 _14026_ (
    .A(_3350__bF$buf3),
    .B(_2_[15]),
    .Y(_3442_)
);

FILL FILL_0__15942_ (
);

FILL FILL_0__15522_ (
);

FILL FILL_0__15102_ (
);

FILL FILL406600x44460 (
);

FILL FILL313880x14820 (
);

FILL FILL500840x79040 (
);

OR2X2 _10786_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .B(_1256__bF$buf4),
    .Y(_1196_)
);

DFFSR _10366_ (
    .CLK(clk_bF$buf112),
    .D(_927_[7]),
    .Q(\datapath_1.regfile_1.regOut[15] [7]),
    .R(rst_bF$buf3),
    .S(vdd)
);

FILL FILL189240x0 (
);

FILL FILL_0__16727_ (
);

FILL FILL_0__16307_ (
);

FILL FILL_0__11862_ (
);

FILL FILL410400x237120 (
);

FILL FILL109440x79040 (
);

FILL FILL235600x291460 (
);

FILL FILL_0__19199_ (
);

OR2X2 _19484_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_8358_)
);

OR2X2 _19064_ (
    .A(_7963_),
    .B(_7956_),
    .Y(_7964_)
);

OR2X2 _8934_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_261_)
);

OR2X2 _8514_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_41_)
);

FILL FILL_1__18519_ (
);

FILL FILL_1__13234_ (
);

XOR2X1 _12932_ (
    .A(_2166_),
    .B(_2369_),
    .Y(_2496_)
);

FILL FILL_0__12227_ (
);

NOR3X1 _12512_ (
    .A(_2101_),
    .B(\control_1.reg_state.dout [1]),
    .C(_2091_),
    .Y(_0_)
);

FILL FILL_1_BUFX2_insert627 (
);

FILL FILL_1_BUFX2_insert629 (
);

DFFSR _9719_ (
    .CLK(clk_bF$buf59),
    .D(_597_[5]),
    .Q(\datapath_1.regfile_1.regOut[10] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL_0__16480_ (
);

AND2X2 _13717_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[18]),
    .Y(_3194_)
);

FILL FILL_1__15800_ (
);

FILL FILL266000x0 (
);

OR2X2 _16189_ (
    .A(_5130_),
    .B(_5131_),
    .Y(_5132_)
);

FILL FILL_1__18272_ (
);

OR2X2 _17970_ (
    .A(_6885_),
    .B(_6886_),
    .Y(_6887_)
);

FILL FILL_0__17265_ (
);

OR2X2 _17550_ (
    .A(_6472_),
    .B(_6471_),
    .Y(_6473_)
);

AND2X2 _17130_ (
    .A(_4223__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_6059_)
);

FILL FILL266760x355680 (
);

OR2X2 _9892_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .B(_794__bF$buf0),
    .Y(_740_)
);

FILL FILL234080x44460 (
);

DFFSR _9472_ (
    .CLK(clk_bF$buf109),
    .D(_465_[16]),
    .Q(\datapath_1.regfile_1.regOut[8] [16]),
    .R(rst_bF$buf84),
    .S(vdd)
);

OR2X2 _9052_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .B(_332__bF$buf2),
    .Y(_320_)
);

FILL FILL166440x19760 (
);

FILL FILL_1__11300_ (
);

OR2X2 _18755_ (
    .A(_7659_),
    .B(_7656_),
    .Y(_7660_)
);

OR2X2 _18335_ (
    .A(_7245_),
    .B(_7242_),
    .Y(_7246_)
);

AND2X2 _13890_ (
    .A(_3326_),
    .B(_3325_),
    .Y(\datapath_1.alu_1.ALUInA [24])
);

FILL FILL_0__13185_ (
);

AND2X2 _13470_ (
    .A(_3002_),
    .B(_2495_),
    .Y(_3003_)
);

OR2X2 _13050_ (
    .A(_2157__bF$buf2),
    .B(_2606_),
    .Y(_2607_)
);

FILL FILL_0__19411_ (
);

FILL FILL117040x83980 (
);

FILL FILL133000x247000 (
);

FILL FILL_1__12925_ (
);

FILL FILL_1__12505_ (
);

FILL FILL_0__9932_ (
);

FILL FILL41800x158080 (
);

FILL FILL47120x232180 (
);

OR2X2 _14675_ (
    .A(vdd),
    .B(\datapath_1.a [16]),
    .Y(_3836_)
);

FILL FILL445360x44460 (
);

OR2X2 _14255_ (
    .A(vdd),
    .B(ALUOut[5]),
    .Y(_3616_)
);

FILL FILL319200x355680 (
);

FILL FILL_0__15751_ (
);

FILL FILL250800x350740 (
);

FILL FILL124640x49400 (
);

AND2X2 _10595_ (
    .A(_1108_),
    .B(_1107_),
    .Y(_1059_[24])
);

AND2X2 _10175_ (
    .A(_888_),
    .B(_887_),
    .Y(_861_[13])
);

FILL FILL_1__17123_ (
);

FILL FILL_0__16956_ (
);

OR2X2 _16821_ (
    .A(_5753_),
    .B(_5754_),
    .Y(_5755_)
);

AND2X2 _16401_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_5341_)
);

FILL FILL_0__16116_ (
);

FILL FILL167200x266760 (
);

FILL FILL254600x271700 (
);

OR2X2 _19293_ (
    .A(_8158_),
    .B(_8189_),
    .Y(_8190_)
);

OR2X2 _8743_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .B(_200__bF$buf4),
    .Y(_154_)
);

FILL FILL264480x217360 (
);

FILL FILL399760x29640 (
);

FILL FILL_1__13883_ (
);

AND2X2 _17606_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_6528_)
);

FILL FILL_0__12876_ (
);

NAND2X1 _12741_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .B(_2272_),
    .Y(_2306_)
);

FILL FILL_0__12456_ (
);

DFFSR _12321_ (
    .CLK(clk_bF$buf104),
    .D(_1917_[27]),
    .Q(\datapath_1.regfile_1.regOut[30] [27]),
    .R(rst_bF$buf80),
    .S(vdd)
);

FILL FILL335920x49400 (
);

FILL FILL49400x187720 (
);

OR2X2 _9948_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_777_)
);

OR2X2 _9528_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_557_)
);

OR2X2 _9108_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_337_)
);

FILL FILL_1__8485_ (
);

FILL FILL128440x49400 (
);

FILL FILL_1__14248_ (
);

FILL FILL_0_BUFX2_insert280 (
);

FILL FILL_0_BUFX2_insert281 (
);

FILL FILL_0_BUFX2_insert282 (
);

FILL FILL459040x172900 (
);

FILL FILL_0_BUFX2_insert284 (
);

AND2X2 _13946_ (
    .A(_3344__bF$buf3),
    .B(gnd),
    .Y(_3373_)
);

OR2X2 _13526_ (
    .A(ALUOut[12]),
    .B(_3079__bF$buf0),
    .Y(_3039_)
);

NOR3X1 _13106_ (
    .A(_2659_),
    .B(_2656_),
    .C(_2657_),
    .Y(_2660_)
);

FILL FILL_0_BUFX2_insert286 (
);

FILL FILL_0_BUFX2_insert288 (
);

FILL FILL231040x202540 (
);

FILL FILL_0__17494_ (
);

FILL FILL_0__17074_ (
);

FILL FILL148200x212420 (
);

FILL FILL_1__16814_ (
);

AND2X2 _9281_ (
    .A(_432_),
    .B(_431_),
    .Y(_399_[16])
);

FILL FILL142120x365560 (
);

FILL FILL_0__15807_ (
);

FILL FILL_0__10522_ (
);

FILL FILL_0__18699_ (
);

OR2X2 _18984_ (
    .A(_7881_),
    .B(_7884_),
    .Y(_7885_)
);

OR2X2 _18564_ (
    .A(_7470_),
    .B(_7471_),
    .Y(_7472_)
);

FILL FILL_0__18279_ (
);

OR2X2 _18144_ (
    .A(_7056_),
    .B(_7057_),
    .Y(_7058_)
);

FILL FILL220400x345800 (
);

FILL FILL156560x326040 (
);

FILL FILL366320x202540 (
);

FILL FILL_0__11727_ (
);

FILL FILL_0__9321_ (
);

FILL FILL_0__11307_ (
);

FILL FILL392160x143260 (
);

FILL FILL60800x138320 (
);

AND2X2 _19349_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_8245_)
);

FILL FILL369360x4940 (
);

FILL FILL163400x296400 (
);

FILL FILL478040x158080 (
);

FILL FILL_0__14199_ (
);

DFFSR _14484_ (
    .CLK(clk_bF$buf2),
    .D(_3672_[19]),
    .Q(\datapath_1.Data [19]),
    .R(rst_bF$buf26),
    .S(vdd)
);

OR2X2 _14064_ (
    .A(_3474_),
    .B(_3471_),
    .Y(\datapath_1.alu_1.ALUInB [20])
);

FILL FILL_0__15980_ (
);

FILL FILL_0__15560_ (
);

FILL FILL77520x281580 (
);

FILL FILL_0__15140_ (
);

FILL FILL47120x49400 (
);

FILL FILL364040x276640 (
);

OR2X2 _15689_ (
    .A(_4639_),
    .B(_4632_),
    .Y(_4640_)
);

OR2X2 _15269_ (
    .A(_4226_),
    .B(_4224_),
    .Y(_4227_)
);

FILL FILL_1__17772_ (
);

FILL FILL_0__16765_ (
);

OR2X2 _16630_ (
    .A(_5563_),
    .B(_5566_),
    .Y(_5567_)
);

FILL FILL_0__16345_ (
);

AND2X2 _16210_ (
    .A(_4197__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_5153_)
);

FILL FILL152760x4940 (
);

FILL FILL465880x74100 (
);

OR2X2 _8972_ (
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .Y(_331_)
);

AND2X2 _8552_ (
    .A(_66_),
    .B(_65_),
    .Y(_3_[31])
);

FILL FILL_1__18137_ (
);

AND2X2 _11189_ (
    .A(_1404_),
    .B(_1403_),
    .Y(_1389_[7])
);

AND2X2 _17835_ (
    .A(_6229__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_6754_)
);

AND2X2 _17415_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_6340_)
);

FILL FILL304000x74100 (
);

NAND2X1 _12970_ (
    .A(_2360_),
    .B(_2504_),
    .Y(_2532_)
);

FILL FILL_0__12685_ (
);

FILL FILL_0__12265_ (
);

AND2X2 _12550_ (
    .A(_2124_),
    .B(\control_1.op [3]),
    .Y(_2138_)
);

OR2X2 _12130_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .B(_1916__bF$buf0),
    .Y(_1892_)
);

FILL FILL_0__18911_ (
);

FILL FILL427120x316160 (
);

FILL FILL307800x266760 (
);

OR2X2 _9757_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_728__bF$buf1),
    .Y(_670_)
);

DFFSR _9337_ (
    .CLK(clk_bF$buf107),
    .D(_399_[10]),
    .Q(\datapath_1.regfile_1.regOut[7] [10]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL22040x148200 (
);

FILL FILL345040x222300 (
);

AND2X2 _13755_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [23]),
    .Y(_3227_)
);

XOR2X1 _13335_ (
    .A(_2186_),
    .B(_2875_),
    .Y(_2876_)
);

FILL FILL_0__14831_ (
);

FILL FILL_0__14411_ (
);

FILL FILL_1__9499_ (
);

FILL FILL_1__16623_ (
);

DFFSR _9090_ (
    .CLK(clk_bF$buf37),
    .D(_267_[21]),
    .Q(\datapath_1.regfile_1.regOut[5] [21]),
    .R(rst_bF$buf46),
    .S(vdd)
);

AND2X2 _15901_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_4849_)
);

FILL FILL_0__15616_ (
);

FILL FILL_1__19095_ (
);

FILL FILL433200x0 (
);

AND2X2 _18793_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_7697_)
);

FILL FILL_0__18088_ (
);

OR2X2 _18373_ (
    .A(_7280_),
    .B(_7283_),
    .Y(_7284_)
);

FILL FILL75240x330980 (
);

FILL FILL66880x207480 (
);

FILL FILL256880x370500 (
);

FILL FILL373920x167960 (
);

FILL FILL202160x103740 (
);

FILL FILL_0__9970_ (
);

FILL FILL_0__9550_ (
);

FILL FILL_0__11956_ (
);

OR2X2 _11821_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .B(_1784__bF$buf4),
    .Y(_1726_)
);

FILL FILL_0__11116_ (
);

DFFSR _11401_ (
    .CLK(clk_bF$buf107),
    .D(_1455_[10]),
    .Q(\datapath_1.regfile_1.regOut[23] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

FILL FILL475000x83980 (
);

AND2X2 _19158_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_8057_)
);

FILL FILL271320x49400 (
);

AND2X2 _14293_ (
    .A(_3641_),
    .B(_3640_),
    .Y(_3606_[17])
);

FILL FILL497040x138320 (
);

OR2X2 _8608_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_134__bF$buf2),
    .Y(_84_)
);

FILL FILL9880x138320 (
);

FILL FILL_1__13748_ (
);

FILL FILL_1__13328_ (
);

FILL FILL300960x44460 (
);

OR2X2 _12606_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(_2170_),
    .Y(_2171_)
);

FILL FILL130720x276640 (
);

AND2X2 _15498_ (
    .A(_4228__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_4452_)
);

AND2X2 _15078_ (
    .A(_4064_),
    .B(_4029_),
    .Y(\datapath_1.regfile_1.regEn [3])
);

FILL FILL320720x59280 (
);

FILL FILL_1__17161_ (
);

FILL FILL309320x370500 (
);

FILL FILL_0__16994_ (
);

FILL FILL_0__16574_ (
);

FILL FILL354920x113620 (
);

FILL FILL37240x113620 (
);

OR2X2 _8781_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_179_)
);

FILL FILL_1__18786_ (
);

FILL FILL_0__17779_ (
);

AND2X2 _17644_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_6566_)
);

FILL FILL_0__17359_ (
);

OR2X2 _17224_ (
    .A(_6147_),
    .B(_6150_),
    .Y(_6151_)
);

FILL FILL_0__12074_ (
);

FILL FILL_0__18720_ (
);

DFFSR _9986_ (
    .CLK(clk_bF$buf52),
    .D(_729_[14]),
    .Q(\datapath_1.regfile_1.regOut[12] [14]),
    .R(rst_bF$buf0),
    .S(vdd)
);

AND2X2 _9566_ (
    .A(_582_),
    .B(_581_),
    .Y(_531_[25])
);

AND2X2 _9146_ (
    .A(_362_),
    .B(_361_),
    .Y(_333_[14])
);

FILL FILL489440x153140 (
);

FILL FILL324520x59280 (
);

FILL FILL_0__10807_ (
);

FILL FILL_0_BUFX2_insert660 (
);

AND2X2 _18849_ (
    .A(_6317__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_7752_)
);

FILL FILL288800x360620 (
);

FILL FILL_0_BUFX2_insert661 (
);

OR2X2 _18429_ (
    .A(_7336_),
    .B(_7338_),
    .Y(_7339_)
);

FILL FILL_0_BUFX2_insert662 (
);

OR2X2 _18009_ (
    .A(_6921_),
    .B(_6924_),
    .Y(_6925_)
);

AND2X2 _13984_ (
    .A(_3350__bF$buf3),
    .B(_2_[9]),
    .Y(_3406_)
);

FILL FILL_0_BUFX2_insert664 (
);

FILL FILL_0__13699_ (
);

FILL FILL_0__13279_ (
);

OR2X2 _13564_ (
    .A(IorD_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [25]),
    .Y(_3064_)
);

INVX1 _13144_ (
    .A(_2695_),
    .Y(\datapath_1.ALUResult [18])
);

FILL FILL_0_BUFX2_insert666 (
);

FILL FILL_0_BUFX2_insert668 (
);

FILL FILL71440x360620 (
);

FILL FILL269800x197600 (
);

FILL FILL_0__19505_ (
);

FILL FILL_0__14640_ (
);

FILL FILL_0__14220_ (
);

FILL FILL303240x311220 (
);

FILL FILL35720x44460 (
);

OR2X2 _14769_ (
    .A(\datapath_1.rd2 [4]),
    .B(_3935__bF$buf3),
    .Y(_3879_)
);

FILL FILL233320x316160 (
);

DFFSR _14349_ (
    .CLK(clk_bF$buf12),
    .D(_3606_[13]),
    .Q(ALUOut[13]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL320720x321100 (
);

FILL FILL_0__15845_ (
);

FILL FILL_0__15425_ (
);

AND2X2 _15710_ (
    .A(_4183__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_4661_)
);

FILL FILL12160x44460 (
);

FILL FILL_0__10980_ (
);

FILL FILL_0__10560_ (
);

AND2X2 _18182_ (
    .A(_6247__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_7096_)
);

OR2X2 _10689_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_1151_)
);

FILL FILL_1__17637_ (
);

OR2X2 _10269_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_931_)
);

FILL FILL502360x138320 (
);

OR2X2 _16915_ (
    .A(_5846_),
    .B(_5845_),
    .Y(_5847_)
);

FILL FILL246240x128440 (
);

AND2X2 _11630_ (
    .A(_1638_),
    .B(_1637_),
    .Y(_1587_[25])
);

FILL FILL_0__11345_ (
);

AND2X2 _11210_ (
    .A(_1418_),
    .B(_1417_),
    .Y(_1389_[14])
);

OR2X2 _19387_ (
    .A(_8281_),
    .B(_8280_),
    .Y(_8282_)
);

DFFSR _8837_ (
    .CLK(clk_bF$buf32),
    .D(_135_[26]),
    .Q(\datapath_1.regfile_1.regOut[3] [26]),
    .R(rst_bF$buf75),
    .S(vdd)
);

BUFX2 _8417_ (
    .A(_1_[25]),
    .Y(memoryAddress[25])
);

FILL FILL_1__13977_ (
);

FILL FILL_1_CLKBUF1_insert1170 (
);

AND2X2 _12835_ (
    .A(_2395_),
    .B(_2399_),
    .Y(_2400_)
);

OR2X2 _12415_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .B(_2048__bF$buf4),
    .Y(_2042_)
);

FILL FILL286520x222300 (
);

FILL FILL_1_CLKBUF1_insert1178 (
);

FILL FILL103360x143260 (
);

FILL FILL_0__13911_ (
);

FILL FILL_1__17390_ (
);

FILL FILL_0__16383_ (
);

FILL FILL280440x375440 (
);

FILL FILL_1__9940_ (
);

OR2X2 _8590_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .B(_134__bF$buf0),
    .Y(_72_)
);

FILL FILL_1__18595_ (
);

INVX1 _17873_ (
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_6791_)
);

FILL FILL_0__17588_ (
);

AND2X2 _17453_ (
    .A(_6264__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_6378_)
);

FILL FILL_0__17168_ (
);

OR2X2 _17033_ (
    .A(_5962_),
    .B(_5955_),
    .Y(_5963_)
);

FILL FILL98800x148200 (
);

OR2X2 _9795_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_695_)
);

OR2X2 _9375_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_475_)
);

FILL FILL433200x281580 (
);

FILL FILL_1__11203_ (
);

FILL FILL_0__8630_ (
);

FILL FILL_0__10616_ (
);

DFFSR _10901_ (
    .CLK(clk_bF$buf55),
    .D(_1191_[26]),
    .Q(\datapath_1.regfile_1.regOut[19] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

OR2X2 _18658_ (
    .A(_7563_),
    .B(_7562_),
    .Y(_7564_)
);

NOR2X1 _18238_ (
    .A(_6310__bF$buf3),
    .B(_7150_),
    .Y(_7151_)
);

OR2X2 _13793_ (
    .A(_3259_),
    .B(_3256_),
    .Y(\datapath_1.mux_pcsrc.dout [28])
);

AND2X2 _13373_ (
    .A(_2909_),
    .B(_2910_),
    .Y(_2911_)
);

FILL FILL310840x276640 (
);

CLKBUF1 CLKBUF1_insert210 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert211 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert212 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert213 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert214 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert215 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert216 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert217 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert218 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert219 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf4)
);

DFFSR _14998_ (
    .CLK(clk_bF$buf40),
    .D(_3936_[17]),
    .Q(\datapath_1.mux_iord.din0 [17]),
    .R(rst_bF$buf53),
    .S(vdd)
);

AND2X2 _14578_ (
    .A(_3791_),
    .B(_3790_),
    .Y(_3738_[26])
);

OR2X2 _14158_ (
    .A(MemToReg_bF$buf4),
    .B(ALUOut[5]),
    .Y(_3550_)
);

FILL FILL227240x54340 (
);

FILL FILL_1__16241_ (
);

FILL FILL159600x29640 (
);

FILL FILL_0__15234_ (
);

DFFSR _10498_ (
    .CLK(clk_bF$buf33),
    .D(_993_[10]),
    .Q(\datapath_1.regfile_1.regOut[16] [10]),
    .R(rst_bF$buf66),
    .S(vdd)
);

OR2X2 _10078_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_860__bF$buf4),
    .Y(_844_)
);

FILL FILL_0__16859_ (
);

FILL FILL_0__16439_ (
);

AND2X2 _16724_ (
    .A(_4187__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_5659_)
);

AND2X2 _16304_ (
    .A(_4217__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_5246_)
);

AND2X2 _19196_ (
    .A(_6259__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_8094_)
);

FILL FILL_0__17800_ (
);

OR2X2 _8646_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_109_)
);

FILL FILL_1__13366_ (
);

OR2X2 _17929_ (
    .A(_6813_),
    .B(_6846_),
    .Y(_6847_)
);

OR2X2 _17509_ (
    .A(_6431_),
    .B(_6432_),
    .Y(_6433_)
);

AND2X2 _12644_ (
    .A(_2201_),
    .B(_2208_),
    .Y(_2209_)
);

FILL FILL_0__12359_ (
);

AND2X2 _12224_ (
    .A(_1934_),
    .B(_1933_),
    .Y(_1917_[8])
);

FILL FILL_0__13720_ (
);

FILL FILL_0__13300_ (
);

FILL FILL_0_BUFX2_insert1011 (
);

FILL FILL_0__16192_ (
);

FILL FILL_0_BUFX2_insert1013 (
);

FILL FILL_0_BUFX2_insert1014 (
);

FILL FILL_0_BUFX2_insert1015 (
);

FILL FILL_0_BUFX2_insert1016 (
);

FILL FILL_0_BUFX2_insert1017 (
);

FILL FILL_0_BUFX2_insert1019 (
);

OR2X2 _13849_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [11]),
    .Y(_3299_)
);

INVX1 _13429_ (
    .A(_2963_),
    .Y(\datapath_1.ALUResult [1])
);

OR2X2 _13009_ (
    .A(_2387__bF$buf2),
    .B(_2568_),
    .Y(_2569_)
);

FILL FILL_0__14925_ (
);

FILL FILL183920x207480 (
);

FILL FILL_0__17397_ (
);

NOR2X1 _17682_ (
    .A(_6310__bF$buf4),
    .B(_6602_),
    .Y(_6603_)
);

FILL FILL36480x74100 (
);

OR2X2 _17262_ (
    .A(_6187_),
    .B(_6188_),
    .Y(_6189_)
);

FILL FILL452960x163020 (
);

FILL FILL257640x123500 (
);

OR2X2 _9184_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .B(_398__bF$buf3),
    .Y(_388_)
);

FILL FILL443840x138320 (
);

FILL FILL187720x128440 (
);

FILL FILL_0__10845_ (
);

OR2X2 _10710_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_1165_)
);

FILL FILL_0__10425_ (
);

FILL FILL_0__10005_ (
);

INVX1 _18887_ (
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_7790_)
);

AND2X2 _18467_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_7376_)
);

OR2X2 _18047_ (
    .A(_6962_),
    .B(_6961_),
    .Y(_6963_)
);

OR2X2 _13182_ (
    .A(_2216_),
    .B(_2730_),
    .Y(_2731_)
);

FILL FILL289560x54340 (
);

FILL FILL_0__19123_ (
);

FILL FILL255360x197600 (
);

DFFSR _11915_ (
    .CLK(clk_bF$buf52),
    .D(_1719_[8]),
    .Q(\datapath_1.regfile_1.regOut[27] [8]),
    .R(rst_bF$buf1),
    .S(vdd)
);

OR2X2 _14387_ (
    .A(vdd),
    .B(\datapath_1.Data [6]),
    .Y(_3684_)
);

FILL FILL505400x163020 (
);

FILL FILL_1__16890_ (
);

FILL FILL_0__15463_ (
);

FILL FILL57760x98800 (
);

FILL FILL418760x143260 (
);

FILL FILL_1__17255_ (
);

FILL FILL269800x24700 (
);

FILL FILL_0__16668_ (
);

OR2X2 _16953_ (
    .A(_5853_),
    .B(_5884_),
    .Y(_5885_)
);

AND2X2 _16533_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_5471_)
);

FILL FILL_0__16248_ (
);

FILL FILL262960x133380 (
);

AND2X2 _16113_ (
    .A(_4210__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_5058_)
);

OR2X2 _8875_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_266__bF$buf3),
    .Y(_222_)
);

BUFX2 _8455_ (
    .A(_2_[31]),
    .Y(memoryWriteData[31])
);

OR2X2 _17738_ (
    .A(_6657_),
    .B(_6656_),
    .Y(_6658_)
);

AND2X2 _17318_ (
    .A(_6243_),
    .B(_6201_),
    .Y(_6244_)
);

FILL FILL_0__12588_ (
);

AND2X2 _12873_ (
    .A(_2437_),
    .B(_2435_),
    .Y(_2438_)
);

FILL FILL_1__19401_ (
);

DFFSR _12453_ (
    .CLK(clk_bF$buf108),
    .D(_1983_[30]),
    .Q(\datapath_1.regfile_1.regOut[31] [30]),
    .R(rst_bF$buf93),
    .S(vdd)
);

OR2X2 _12033_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_1847_)
);

FILL FILL430920x98800 (
);

FILL FILL272080x222300 (
);

FILL FILL_0__8915_ (
);

AND2X2 _13658_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3144_)
);

NOR2X1 _13238_ (
    .A(_2764_),
    .B(_2498_),
    .Y(_2784_)
);

FILL FILL_1__15741_ (
);

FILL FILL_0__14314_ (
);

FILL FILL452960x256880 (
);

OR2X2 _17491_ (
    .A(_6406_),
    .B(_6414_),
    .Y(_6415_)
);

OR2X2 _17071_ (
    .A(_6000_),
    .B(_5997_),
    .Y(_6001_)
);

FILL FILL439280x167960 (
);

FILL FILL201400x251940 (
);

FILL FILL_1__16106_ (
);

FILL FILL_0__15939_ (
);

AND2X2 _15804_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_4753_)
);

FILL FILL_0__10654_ (
);

AND2X2 _18696_ (
    .A(_6262__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_7602_)
);

AND2X2 _18276_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_7188_)
);

FILL FILL_0__19352_ (
);

FILL FILL_1__12866_ (
);

FILL FILL262200x9880 (
);

FILL FILL505400x256880 (
);

FILL FILL_0__9453_ (
);

FILL FILL_0__11859_ (
);

FILL FILL141360x247000 (
);

FILL FILL171760x158080 (
);

FILL FILL_0__9033_ (
);

OR2X2 _11724_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_1681_)
);

FILL FILL_0__11439_ (
);

FILL FILL456000x301340 (
);

OR2X2 _11304_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_1461_)
);

AND2X2 _14196_ (
    .A(_3575_),
    .B(_3574_),
    .Y(\datapath_1.mux_wd3.dout [17])
);

FILL FILL437000x138320 (
);

FILL FILL146680x34580 (
);

FILL FILL_0__15692_ (
);

FILL FILL_1_BUFX2_insert590 (
);

FILL FILL72960x242060 (
);

FILL FILL_1_BUFX2_insert592 (
);

AND2X2 _12929_ (
    .A(_2493_),
    .B(_2385_),
    .Y(_2494_)
);

INVX2 _12509_ (
    .A(_2104_),
    .Y(MemToReg)
);

FILL FILL_1_BUFX2_insert594 (
);

FILL FILL249280x0 (
);

FILL FILL376960x153140 (
);

FILL FILL_0__16897_ (
);

AND2X2 _16762_ (
    .A(_5696_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [23])
);

FILL FILL_0__16057_ (
);

OR2X2 _16342_ (
    .A(_5282_),
    .B(_5281_),
    .Y(_5283_)
);

FILL FILL281960x113620 (
);

DFFSR _8684_ (
    .CLK(clk_bF$buf111),
    .D(_69_[2]),
    .Q(\datapath_1.regfile_1.regOut[2] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

FILL FILL348840x286520 (
);

FILL FILL_1__18689_ (
);

BUFX2 BUFX2_insert260 (
    .A(_6271_),
    .Y(_6271__bF$buf3)
);

BUFX2 BUFX2_insert261 (
    .A(_6271_),
    .Y(_6271__bF$buf2)
);

BUFX2 BUFX2_insert262 (
    .A(_6271_),
    .Y(_6271__bF$buf1)
);

BUFX2 BUFX2_insert263 (
    .A(_6271_),
    .Y(_6271__bF$buf0)
);

BUFX2 BUFX2_insert264 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf4 )
);

OR2X2 _17967_ (
    .A(_6880_),
    .B(_6883_),
    .Y(_6884_)
);

OR2X2 _17547_ (
    .A(_6466_),
    .B(_6469_),
    .Y(_6470_)
);

BUFX2 BUFX2_insert265 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf3 )
);

BUFX2 BUFX2_insert266 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf2 )
);

OR2X2 _17127_ (
    .A(_6052_),
    .B(_6055_),
    .Y(_6056_)
);

BUFX2 BUFX2_insert267 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf1 )
);

FILL FILL198360x350740 (
);

FILL FILL120840x316160 (
);

BUFX2 BUFX2_insert268 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf0 )
);

BUFX2 BUFX2_insert269 (
    .A(_2379_),
    .Y(_2379__bF$buf3)
);

INVX1 _12682_ (
    .A(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2247_)
);

FILL FILL297160x0 (
);

OR2X2 _12262_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .B(_1982__bF$buf0),
    .Y(_1960_)
);

FILL FILL_0__18623_ (
);

FILL FILL_0__18203_ (
);

FILL FILL179360x187720 (
);

FILL FILL330600x19760 (
);

FILL FILL384560x365560 (
);

FILL FILL256120x133380 (
);

OR2X2 _9889_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .B(_794__bF$buf4),
    .Y(_738_)
);

DFFSR _9469_ (
    .CLK(clk_bF$buf61),
    .D(_465_[13]),
    .Q(\datapath_1.regfile_1.regOut[8] [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

OR2X2 _9049_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .B(_332__bF$buf0),
    .Y(_318_)
);

FILL FILL_0__8724_ (
);

FILL FILL_1__14189_ (
);

AND2X2 _13887_ (
    .A(_3324_),
    .B(_3323_),
    .Y(\datapath_1.alu_1.ALUInA [23])
);

AND2X2 _13467_ (
    .A(_2999_),
    .B(_2983_),
    .Y(_3000_)
);

OR2X2 _13047_ (
    .A(_2264_),
    .B(_2603_),
    .Y(_2604_)
);

FILL FILL_0__19408_ (
);

FILL FILL_0__14963_ (
);

FILL FILL_0__14543_ (
);

FILL FILL_0__9509_ (
);

FILL FILL412680x222300 (
);

FILL FILL_1__16755_ (
);

FILL FILL_1__11890_ (
);

FILL FILL342760x227240 (
);

FILL FILL_0__15328_ (
);

OR2X2 _15613_ (
    .A(_4563_),
    .B(_4564_),
    .Y(_4565_)
);

FILL FILL334400x19760 (
);

FILL FILL_0__10043_ (
);

AND2X2 _18085_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_7000_)
);

FILL FILL_0__19161_ (
);

FILL FILL173280x128440 (
);

FILL FILL102600x291460 (
);

FILL FILL_1__12255_ (
);

FILL FILL254600x34580 (
);

OR2X2 _16818_ (
    .A(_5751_),
    .B(_5750_),
    .Y(_5752_)
);

FILL FILL_0__9682_ (
);

FILL FILL_1__18901_ (
);

OR2X2 _11953_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .B(_1850__bF$buf3),
    .Y(_1794_)
);

DFFSR _11533_ (
    .CLK(clk_bF$buf34),
    .D(_1521_[13]),
    .Q(\datapath_1.regfile_1.regOut[24] [13]),
    .R(rst_bF$buf70),
    .S(vdd)
);

FILL FILL_0__11248_ (
);

OR2X2 _11113_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_1388__bF$buf4),
    .Y(_1374_)
);

FILL FILL190760x138320 (
);

FILL FILL429400x44460 (
);

FILL FILL164920x69160 (
);

FILL FILL294120x167960 (
);

FILL FILL_0__15081_ (
);

OR2X2 _12738_ (
    .A(_2276_),
    .B(_2302_),
    .Y(_2303_)
);

DFFSR _12318_ (
    .CLK(clk_bF$buf35),
    .D(_1917_[24]),
    .Q(\datapath_1.regfile_1.regOut[30] [24]),
    .R(rst_bF$buf67),
    .S(vdd)
);

FILL FILL_1__14401_ (
);

FILL FILL317680x232180 (
);

FILL FILL_0__13814_ (
);

OR2X2 _16991_ (
    .A(_5921_),
    .B(_5920_),
    .Y(_5922_)
);

AND2X2 _16571_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_5508_)
);

FILL FILL_0__16286_ (
);

OR2X2 _16151_ (
    .A(_5094_),
    .B(_5091_),
    .Y(_5095_)
);

FILL FILL_1__9003_ (
);

OR2X2 _8493_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_27_)
);

FILL FILL_1__15606_ (
);

FILL FILL203680x350740 (
);

FILL FILL_1__18078_ (
);

OR2X2 _17776_ (
    .A(_6694_),
    .B(_6695_),
    .Y(_6696_)
);

AND2X2 _17356_ (
    .A(_6274_),
    .B(_6281_),
    .Y(_6282_)
);

NOR2X1 _12491_ (
    .A(_2094_),
    .B(\control_1.reg_state.dout [0]),
    .Y(Branch)
);

AND2X2 _12071_ (
    .A(_1852_),
    .B(_1915_),
    .Y(_1851_[0])
);

FILL FILL_0__18852_ (
);

FILL FILL_0__18012_ (
);

AND2X2 _9698_ (
    .A(_650_),
    .B(_649_),
    .Y(_597_[26])
);

AND2X2 _9278_ (
    .A(_430_),
    .B(_429_),
    .Y(_399_[15])
);

FILL FILL_1__11946_ (
);

FILL FILL_0__10939_ (
);

OR2X2 _10804_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .B(_1256__bF$buf3),
    .Y(_1208_)
);

AND2X2 _13696_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[15]),
    .Y(_3176_)
);

INVX1 _13276_ (
    .A(_2819_),
    .Y(\datapath_1.ALUResult [10])
);

FILL FILL63840x54340 (
);

FILL FILL338960x350740 (
);

FILL FILL60800x251940 (
);

FILL FILL_0__19217_ (
);

OR2X2 _19502_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [25]),
    .Y(_8370_)
);

FILL FILL_0__14772_ (
);

FILL FILL114000x316160 (
);

FILL FILL319960x187720 (
);

FILL FILL_0__9318_ (
);

FILL FILL100320x340860 (
);

FILL FILL456760x247000 (
);

FILL FILL_0__15977_ (
);

AND2X2 _15842_ (
    .A(_4210__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_4791_)
);

FILL FILL_0__15557_ (
);

AND2X2 _15422_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_4377_)
);

DFFSR _15002_ (
    .CLK(clk_bF$buf77),
    .D(_3936_[21]),
    .Q(\datapath_1.mux_iord.din0 [21]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__10692_ (
);

FILL FILL290320x197600 (
);

FILL FILL120080x49400 (
);

FILL FILL49400x232180 (
);

AND2X2 _16627_ (
    .A(_4230__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_5564_)
);

OR2X2 _16207_ (
    .A(_5148_),
    .B(_5149_),
    .Y(_5150_)
);

FILL FILL_0__11897_ (
);

FILL FILL_0__9491_ (
);

AND2X2 _11762_ (
    .A(_1706_),
    .B(_1705_),
    .Y(_1653_[26])
);

FILL FILL_0__11477_ (
);

AND2X2 _11342_ (
    .A(_1486_),
    .B(_1485_),
    .Y(_1455_[15])
);

FILL FILL_0__11057_ (
);

OR2X2 _19099_ (
    .A(_7965_),
    .B(_7998_),
    .Y(_7999_)
);

FILL FILL_0__17703_ (
);

DFFSR _8969_ (
    .CLK(clk_bF$buf64),
    .D(_201_[29]),
    .Q(\datapath_1.regfile_1.regOut[4] [29]),
    .R(rst_bF$buf73),
    .S(vdd)
);

AND2X2 _8549_ (
    .A(_64_),
    .B(_63_),
    .Y(_3_[30])
);

OR2X2 _9910_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .B(_794__bF$buf4),
    .Y(_752_)
);

FILL FILL313880x128440 (
);

FILL FILL_1_BUFX2_insert970 (
);

XOR2X1 _12967_ (
    .A(_2359_),
    .B(_2350_),
    .Y(_2529_)
);

FILL FILL_1_BUFX2_insert972 (
);

AND2X2 _12547_ (
    .A(_2135_),
    .B(_2118_),
    .Y(_2136_)
);

OR2X2 _12127_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .B(_1916__bF$buf4),
    .Y(_1890_)
);

FILL FILL_1_BUFX2_insert974 (
);

FILL FILL252320x256880 (
);

FILL FILL_1__14210_ (
);

FILL FILL_0__13203_ (
);

AND2X2 _16380_ (
    .A(_4239__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_5320_)
);

FILL FILL266760x217360 (
);

FILL FILL214320x88920 (
);

FILL FILL_1__15835_ (
);

FILL FILL_1__10970_ (
);

FILL FILL_0__14408_ (
);

BUFX2 BUFX2_insert640 (
    .A(_6244_),
    .Y(_6244__bF$buf4)
);

BUFX2 BUFX2_insert641 (
    .A(_6244_),
    .Y(_6244__bF$buf3)
);

BUFX2 BUFX2_insert642 (
    .A(_6244_),
    .Y(_6244__bF$buf2)
);

BUFX2 BUFX2_insert643 (
    .A(_6244_),
    .Y(_6244__bF$buf1)
);

BUFX2 BUFX2_insert644 (
    .A(_6244_),
    .Y(_6244__bF$buf0)
);

BUFX2 BUFX2_insert645 (
    .A(_6282_),
    .Y(_6282__bF$buf4)
);

OR2X2 _17585_ (
    .A(_6507_),
    .B(_6504_),
    .Y(_6508_)
);

BUFX2 BUFX2_insert646 (
    .A(_6282_),
    .Y(_6282__bF$buf3)
);

AND2X2 _17165_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_6093_)
);

BUFX2 BUFX2_insert647 (
    .A(_6282_),
    .Y(_6282__bF$buf2)
);

BUFX2 BUFX2_insert648 (
    .A(_6282_),
    .Y(_6282__bF$buf1)
);

BUFX2 BUFX2_insert649 (
    .A(_6282_),
    .Y(_6282__bF$buf0)
);

FILL FILL_0__18661_ (
);

FILL FILL277400x0 (
);

FILL FILL_0__18241_ (
);

FILL FILL402800x301340 (
);

DFFSR _9087_ (
    .CLK(clk_bF$buf67),
    .D(_267_[18]),
    .Q(\datapath_1.regfile_1.regOut[5] [18]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_1__11335_ (
);

FILL FILL_0__8762_ (
);

FILL FILL_0__10328_ (
);

AND2X2 _10613_ (
    .A(_1120_),
    .B(_1119_),
    .Y(_1059_[30])
);

FILL FILL402040x207480 (
);

FILL FILL172520x232180 (
);

NAND2X1 _13085_ (
    .A(_2466_),
    .B(_2548_),
    .Y(_2640_)
);

FILL FILL_0__19446_ (
);

FILL FILL218120x88920 (
);

FILL FILL_0__19026_ (
);

OR2X2 _19311_ (
    .A(_8199_),
    .B(_8206_),
    .Y(_8207_)
);

FILL FILL491720x177840 (
);

FILL FILL482600x79040 (
);

FILL FILL_0__14161_ (
);

FILL FILL_0__9967_ (
);

FILL FILL_0__9127_ (
);

OR2X2 _11818_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .B(_1784__bF$buf4),
    .Y(_1724_)
);

FILL FILL144400x365560 (
);

FILL FILL231800x370500 (
);

FILL FILL345800x118560 (
);

FILL FILL_0__15786_ (
);

FILL FILL_0__15366_ (
);

OR2X2 _15651_ (
    .A(_4602_),
    .B(_4601_),
    .Y(_4603_)
);

NOR3X1 _15231_ (
    .A(_4144_),
    .B(_4140_),
    .C(_4153_),
    .Y(_4189_)
);

FILL FILL231040x276640 (
);

FILL FILL3800x301340 (
);

FILL FILL82840x24700 (
);

FILL FILL368600x202540 (
);

FILL FILL_1__17578_ (
);

OR2X2 _16856_ (
    .A(_5788_),
    .B(_5781_),
    .Y(_5789_)
);

FILL FILL68400x212420 (
);

AND2X2 _16436_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_5376_)
);

OR2X2 _16016_ (
    .A(_4961_),
    .B(_4958_),
    .Y(_4962_)
);

FILL FILL486400x79040 (
);

FILL FILL199120x103740 (
);

OR2X2 _11991_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_1819_)
);

OR2X2 _11571_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_1599_)
);

FILL FILL81320x207480 (
);

DFFSR _11151_ (
    .CLK(clk_bF$buf3),
    .D(_1323_[18]),
    .Q(\datapath_1.regfile_1.regOut[21] [18]),
    .R(rst_bF$buf4),
    .S(vdd)
);

FILL FILL79800x281580 (
);

OR2X2 _8778_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_177_)
);

FILL FILL_1__10606_ (
);

NAND2X1 _12776_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(_2340_),
    .Y(_2341_)
);

AND2X2 _12356_ (
    .A(_2002_),
    .B(_2001_),
    .Y(_1983_[9])
);

FILL FILL_0__18717_ (
);

FILL FILL_0__13852_ (
);

FILL FILL383800x286520 (
);

FILL FILL_0__13432_ (
);

FILL FILL66120x286520 (
);

FILL FILL_1__15224_ (
);

OR2X2 _14922_ (
    .A(\datapath_1.mux_pcsrc.dout [12]),
    .B(_4001__bF$buf3),
    .Y(_3961_)
);

FILL FILL_0__14217_ (
);

OR2X2 _14502_ (
    .A(memoryOutData[1]),
    .B(_3803__bF$buf0),
    .Y(_3741_)
);

OR2X2 _17394_ (
    .A(_6319_),
    .B(_6314_),
    .Y(_6320_)
);

FILL FILL_0__18890_ (
);

FILL FILL_0__18470_ (
);

FILL FILL_0__18050_ (
);

FILL FILL43320x311220 (
);

FILL FILL24320x148200 (
);

AND2X2 _15707_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_4658_)
);

FILL FILL347320x222300 (
);

FILL FILL_0__8991_ (
);

FILL FILL_0__10977_ (
);

OR2X2 _10842_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_1233_)
);

FILL FILL_0__10557_ (
);

FILL FILL_0__10137_ (
);

OR2X2 _10422_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_1013_)
);

FILL FILL360240x217360 (
);

DFFSR _10002_ (
    .CLK(clk_bF$buf108),
    .D(_729_[30]),
    .Q(\datapath_1.regfile_1.regOut[12] [30]),
    .R(rst_bF$buf93),
    .S(vdd)
);

AND2X2 _18599_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_7506_)
);

NOR2X1 _18179_ (
    .A(_6310__bF$buf2),
    .B(_7092_),
    .Y(_7093_)
);

FILL FILL237880x118560 (
);

DFFSR _19540_ (
    .CLK(clk_bF$buf65),
    .D(_8320_[17]),
    .Q(\datapath_1.regfile_1.regOut[0] [17]),
    .R(rst_bF$buf31),
    .S(vdd)
);

OR2X2 _19120_ (
    .A(_8015_),
    .B(_8018_),
    .Y(_8019_)
);

FILL FILL60040x227240 (
);

FILL FILL_1__12349_ (
);

FILL FILL_0__9776_ (
);

FILL FILL111720x158080 (
);

AND2X2 _11627_ (
    .A(_1636_),
    .B(_1635_),
    .Y(_1587_[24])
);

AND2X2 _11207_ (
    .A(_1416_),
    .B(_1415_),
    .Y(_1389_[13])
);

FILL FILL163400x345800 (
);

OR2X2 _14099_ (
    .A(_3504_),
    .B(_3501_),
    .Y(\datapath_1.alu_1.ALUInB [25])
);

FILL FILL_0__12703_ (
);

FILL FILL_1__16182_ (
);

OR2X2 _15880_ (
    .A(_4824_),
    .B(_4827_),
    .Y(_4828_)
);

FILL FILL66880x19760 (
);

AND2X2 _15460_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_4415_)
);

FILL FILL_0__15175_ (
);

FILL FILL77520x330980 (
);

AND2X2 _15040_ (
    .A(_4016_),
    .B(_4028_),
    .Y(_4029_)
);

FILL FILL17480x83980 (
);

OR2X2 _16665_ (
    .A(_5600_),
    .B(_5585_),
    .Y(_5601_)
);

FILL FILL324520x9880 (
);

OR2X2 _16245_ (
    .A(_5187_),
    .B(_5186_),
    .Y(_5188_)
);

FILL FILL294120x49400 (
);

FILL FILL499320x138320 (
);

OR2X2 _11380_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .B(_1520__bF$buf4),
    .Y(_1512_)
);

FILL FILL_0__11095_ (
);

FILL FILL307800x128440 (
);

FILL FILL_0__17741_ (
);

FILL FILL_0__17321_ (
);

FILL FILL304000x9880 (
);

OR2X2 _8587_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(_134__bF$buf0),
    .Y(_70_)
);

FILL FILL_1__10415_ (
);

FILL FILL343520x59280 (
);

DFFSR _12585_ (
    .CLK(clk_bF$buf20),
    .D(_2143_[1]),
    .Q(\control_1.reg_state.dout [1]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _12165_ (
    .CLK(clk_bF$buf41),
    .D(_1851_[0]),
    .Q(\datapath_1.regfile_1.regOut[29] [0]),
    .R(rst_bF$buf63),
    .S(vdd)
);

FILL FILL_0__18946_ (
);

FILL FILL339720x103740 (
);

AND2X2 _18811_ (
    .A(_6232__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_7715_)
);

FILL FILL_0__18526_ (
);

FILL FILL206720x83980 (
);

FILL FILL_1__9690_ (
);

FILL FILL52440x108680 (
);

FILL FILL326800x4940 (
);

FILL FILL_1__15873_ (
);

DFFSR _14731_ (
    .CLK(clk_bF$buf38),
    .D(_3804_[8]),
    .Q(\datapath_1.a [8]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL_0__14446_ (
);

FILL FILL_0__14026_ (
);

AND2X2 _14311_ (
    .A(_3653_),
    .B(_3652_),
    .Y(_3606_[23])
);

CLKBUF1 CLKBUF1_insert180 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert181 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert182 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert183 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert184 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert185 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf38)
);

FILL FILL31160x44460 (
);

CLKBUF1 CLKBUF1_insert186 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert187 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert188 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert189 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf34)
);

FILL FILL347320x59280 (
);

OR2X2 _15936_ (
    .A(_4881_),
    .B(_4882_),
    .Y(_4883_)
);

OR2X2 _15516_ (
    .A(_4468_),
    .B(_4469_),
    .Y(_4470_)
);

FILL FILL_0__10786_ (
);

OR2X2 _10651_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(_1190__bF$buf1),
    .Y(_1126_)
);

DFFSR _10231_ (
    .CLK(clk_bF$buf28),
    .D(_861_[1]),
    .Q(\datapath_1.regfile_1.regOut[14] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL491720x247000 (
);

FILL FILL_0__19064_ (
);

FILL FILL113240x128440 (
);

FILL FILL_1__12578_ (
);

FILL FILL_0__9165_ (
);

OR2X2 _11856_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[27] [15]),
    .Y(_1749_)
);

OR2X2 _11436_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_1529_)
);

DFFSR _11016_ (
    .CLK(clk_bF$buf113),
    .D(_1257_[12]),
    .Q(\datapath_1.regfile_1.regOut[20] [12]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_0__12932_ (
);

FILL FILL_0__12512_ (
);

FILL FILL504640x138320 (
);

FILL FILL_0__13717_ (
);

FILL FILL_1__17196_ (
);

AND2X2 _16894_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .Y(_5826_)
);

AND2X2 _16474_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_5413_)
);

OR2X2 _16054_ (
    .A(_4999_),
    .B(_4996_),
    .Y(_5000_)
);

FILL FILL_0__17970_ (
);

FILL FILL_0__17130_ (
);

FILL FILL371640x212420 (
);

BUFX2 _8396_ (
    .A(_1_[4]),
    .Y(memoryAddress[4])
);

FILL FILL198360x59280 (
);

FILL FILL329840x24700 (
);

FILL FILL382280x59280 (
);

FILL FILL_1__10224_ (
);

FILL FILL15200x14820 (
);

FILL FILL288800x222300 (
);

AND2X2 _17679_ (
    .A(_6328__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_6600_)
);

OR2X2 _17259_ (
    .A(_6184_),
    .B(_6185_),
    .Y(_6186_)
);

OR2X2 _12394_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .B(_2048__bF$buf3),
    .Y(_2028_)
);

FILL FILL_1__19342_ (
);

AND2X2 _18620_ (
    .A(_6326__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_7527_)
);

FILL FILL_0__18335_ (
);

OR2X2 _18200_ (
    .A(_7111_),
    .B(_7112_),
    .Y(_7113_)
);

FILL FILL282720x375440 (
);

FILL FILL_0__13470_ (
);

FILL FILL_0__13050_ (
);

FILL FILL_0__8856_ (
);

FILL FILL_0__8436_ (
);

OR2X2 _10707_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_1163_)
);

AND2X2 _13599_ (
    .A(_3084__bF$buf1),
    .B(gnd),
    .Y(_3093_)
);

NAND2X1 _13179_ (
    .A(\datapath_1.alu_1.ALUInA [14]),
    .B(_2252_),
    .Y(_2728_)
);

OR2X2 _19405_ (
    .A(_8296_),
    .B(_8299_),
    .Y(_8300_)
);

OR2X2 _14960_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [25]),
    .Y(_3986_)
);

FILL FILL_0__14675_ (
);

FILL FILL_0__14255_ (
);

OR2X2 _14540_ (
    .A(IRWrite_bF$buf0),
    .B(\datapath_1.PCJump [16]),
    .Y(_3766_)
);

OR2X2 _14120_ (
    .A(_3522_),
    .B(_3519_),
    .Y(\datapath_1.alu_1.ALUInB [28])
);

FILL FILL_1__16047_ (
);

OR2X2 _15745_ (
    .A(_4694_),
    .B(_4691_),
    .Y(_4695_)
);

AND2X2 _15325_ (
    .A(_4230__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_4282_)
);

DFFSR _10880_ (
    .CLK(clk_bF$buf70),
    .D(_1191_[5]),
    .Q(\datapath_1.regfile_1.regOut[19] [5]),
    .R(rst_bF$buf66),
    .S(vdd)
);

AND2X2 _10460_ (
    .A(_1038_),
    .B(_1037_),
    .Y(_993_[22])
);

FILL FILL_0__10175_ (
);

AND2X2 _10040_ (
    .A(_818_),
    .B(_817_),
    .Y(_795_[11])
);

FILL FILL_0__16821_ (
);

FILL FILL263720x321100 (
);

FILL FILL_0__19293_ (
);

FILL FILL_1__12387_ (
);

FILL FILL193800x326040 (
);

DFFSR _11665_ (
    .CLK(clk_bF$buf5),
    .D(_1587_[16]),
    .Q(\datapath_1.regfile_1.regOut[25] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

OR2X2 _11245_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_1454__bF$buf0),
    .Y(_1442_)
);

FILL FILL_0__17606_ (
);

FILL FILL490200x113620 (
);

OR2X2 _9813_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_707_)
);

FILL FILL_1__8770_ (
);

FILL FILL_1__14533_ (
);

FILL FILL348840x172900 (
);

FILL FILL_0__13946_ (
);

AND2X2 _13811_ (
    .A(_3087__bF$buf1),
    .B(\datapath_1.ALUResult [31]),
    .Y(_3275_)
);

FILL FILL_0__13526_ (
);

AND2X2 _16283_ (
    .A(_4223__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_5225_)
);

FILL FILL_1__9135_ (
);

FILL FILL120080x108680 (
);

FILL FILL_1__10033_ (
);

FILL FILL6080x261820 (
);

FILL FILL284240x345800 (
);

AND2X2 _17488_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_6412_)
);

AND2X2 _17068_ (
    .A(_4195__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_5998_)
);

FILL FILL_0__18984_ (
);

FILL FILL_0__18564_ (
);

FILL FILL_0__18144_ (
);

FILL FILL433200x330980 (
);

OR2X2 _10936_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .B(_1322__bF$buf1),
    .Y(_1276_)
);

DFFSR _10516_ (
    .CLK(clk_bF$buf91),
    .D(_993_[28]),
    .Q(\datapath_1.regfile_1.regOut[16] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL310080x365560 (
);

OR2X2 _19214_ (
    .A(_8111_),
    .B(_8109_),
    .Y(_8112_)
);

FILL FILL473480x232180 (
);

FILL FILL259920x123500 (
);

FILL FILL42560x123500 (
);

FILL FILL_1__16696_ (
);

FILL FILL_1__16276_ (
);

OR2X2 _15974_ (
    .A(_4920_),
    .B(_4919_),
    .Y(_4921_)
);

FILL FILL_0__15269_ (
);

AND2X2 _15554_ (
    .A(_4214__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_4507_)
);

NOR2X1 _15134_ (
    .A(_4106_),
    .B(_4042_),
    .Y(\datapath_1.regfile_1.regEn [17])
);

FILL FILL472720x24700 (
);

FILL FILL445360x365560 (
);

FILL FILL_0__16210_ (
);

FILL FILL340480x187720 (
);

FILL FILL265240x24700 (
);

FILL FILL257640x197600 (
);

OR2X2 _16759_ (
    .A(_5686_),
    .B(_5693_),
    .Y(_5694_)
);

OR2X2 _16339_ (
    .A(_5279_),
    .B(_5278_),
    .Y(_5280_)
);

AND2X2 _11894_ (
    .A(_1774_),
    .B(_1773_),
    .Y(_1719_[27])
);

FILL FILL_0__11189_ (
);

AND2X2 _11474_ (
    .A(_1554_),
    .B(_1553_),
    .Y(_1521_[16])
);

AND2X2 _11054_ (
    .A(_1334_),
    .B(_1333_),
    .Y(_1323_[5])
);

FILL FILL_0__17835_ (
);

FILL FILL_0__17415_ (
);

OR2X2 _17700_ (
    .A(_6620_),
    .B(_6607_),
    .Y(_6621_)
);

FILL FILL_0__12970_ (
);

FILL FILL_0__12550_ (
);

OR2X2 _9622_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .B(_662__bF$buf3),
    .Y(_600_)
);

DFFSR _9202_ (
    .CLK(clk_bF$buf79),
    .D(_333_[4]),
    .Q(\datapath_1.regfile_1.regOut[6] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

INVX1 _12679_ (
    .A(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2244_)
);

FILL FILL_1__19207_ (
);

OR2X2 _12259_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_1982__bF$buf4),
    .Y(_1958_)
);

FILL FILL107160x34580 (
);

AND2X2 _18905_ (
    .A(_7807_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd1 [23])
);

FILL FILL147440x217360 (
);

FILL FILL_0__13335_ (
);

AND2X2 _13620_ (
    .A(_3084__bF$buf3),
    .B(\aluControl_1.inst [2]),
    .Y(_3111_)
);

XNOR2X1 _13200_ (
    .A(_2211_),
    .B(_2748_),
    .Y(_2749_)
);

OR2X2 _16092_ (
    .A(_5036_),
    .B(_5035_),
    .Y(_5037_)
);

FILL FILL219640x256880 (
);

FILL FILL57000x103740 (
);

OR2X2 _14825_ (
    .A(vdd),
    .B(_2_[23]),
    .Y(_3916_)
);

OR2X2 _14405_ (
    .A(vdd),
    .B(\datapath_1.Data [12]),
    .Y(_3696_)
);

OR2X2 _17297_ (
    .A(_6217_),
    .B(_6222_),
    .Y(_6223_)
);

FILL FILL268280x281580 (
);

FILL FILL_0__18793_ (
);

FILL FILL274360x222300 (
);

FILL FILL_1__11467_ (
);

FILL FILL245480x19760 (
);

FILL FILL_0__8894_ (
);

AND2X2 _10745_ (
    .A(_1188_),
    .B(_1187_),
    .Y(_1125_[31])
);

AND2X2 _10325_ (
    .A(_968_),
    .B(_967_),
    .Y(_927_[20])
);

FILL FILL_0__19158_ (
);

OR2X2 _19443_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8331_)
);

OR2X2 _19023_ (
    .A(_7923_),
    .B(_7920_),
    .Y(_7924_)
);

FILL FILL_0__14293_ (
);

FILL FILL_0__9259_ (
);

FILL FILL_1__13613_ (
);

OR2X2 _15783_ (
    .A(_4732_),
    .B(_4729_),
    .Y(_4733_)
);

FILL FILL_0__15498_ (
);

AND2X2 _15363_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_4319_)
);

FILL FILL412680x158080 (
);

FILL FILL249280x19760 (
);

FILL FILL143640x247000 (
);

OR2X2 _16988_ (
    .A(_5918_),
    .B(_5917_),
    .Y(_5919_)
);

OR2X2 _16568_ (
    .A(_5505_),
    .B(_5490_),
    .Y(_5506_)
);

AND2X2 _16148_ (
    .A(_4187__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_5092_)
);

DFFSR _11283_ (
    .CLK(clk_bF$buf85),
    .D(_1389_[21]),
    .Q(\datapath_1.regfile_1.regOut[22] [21]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL_0__17644_ (
);

FILL FILL_1__10318_ (
);

FILL FILL105640x54340 (
);

DFFSR _9851_ (
    .CLK(clk_bF$buf3),
    .D(_663_[8]),
    .Q(\datapath_1.regfile_1.regOut[11] [8]),
    .R(rst_bF$buf58),
    .S(vdd)
);

AND2X2 _9431_ (
    .A(_512_),
    .B(_511_),
    .Y(_465_[23])
);

AND2X2 _9011_ (
    .A(_292_),
    .B(_291_),
    .Y(_267_[12])
);

FILL FILL_1__19436_ (
);

INVX1 _12488_ (
    .A(\control_1.reg_state.dout [2]),
    .Y(_2093_)
);

OR2X2 _12068_ (
    .A(\datapath_1.regfile_1.regOut[29] [0]),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .Y(_1915_)
);

FILL FILL_1__14571_ (
);

INVX1 _18714_ (
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_7619_)
);

FILL FILL_0__18429_ (
);

FILL FILL_0__18009_ (
);

FILL FILL_0__13984_ (
);

FILL FILL_0__13564_ (
);

FILL FILL_0__13144_ (
);

FILL FILL361000x335920 (
);

FILL FILL433960x276640 (
);

OR2X2 _14634_ (
    .A(\datapath_1.rd1 [2]),
    .B(_3869__bF$buf4),
    .Y(_3809_)
);

AND2X2 _14214_ (
    .A(_3587_),
    .B(_3586_),
    .Y(\datapath_1.mux_wd3.dout [23])
);

FILL FILL_0__15710_ (
);

FILL FILL_0__18182_ (
);

OR2X2 _15839_ (
    .A(_4787_),
    .B(_4786_),
    .Y(_4788_)
);

AND2X2 _15419_ (
    .A(_4200__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_4374_)
);

FILL FILL418760x49400 (
);

OR2X2 _10974_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_1301_)
);

FILL FILL_0__10689_ (
);

OR2X2 _10554_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_1081_)
);

FILL FILL_1__17502_ (
);

FILL FILL_0__10269_ (
);

INVX2 _10134_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .Y(_926_)
);

FILL FILL_0__11630_ (
);

FILL FILL_0__11210_ (
);

FILL FILL_0__19387_ (
);

INVX1 _19252_ (
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_8149_)
);

FILL FILL250040x34580 (
);

DFFSR _8702_ (
    .CLK(clk_bF$buf10),
    .D(_69_[20]),
    .Q(\datapath_1.regfile_1.regOut[2] [20]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL414960x222300 (
);

AND2X2 _11759_ (
    .A(_1704_),
    .B(_1703_),
    .Y(_1653_[25])
);

AND2X2 _11339_ (
    .A(_1484_),
    .B(_1483_),
    .Y(_1455_[14])
);

FILL FILL_1__13842_ (
);

FILL FILL30400x276640 (
);

FILL FILL27360x227240 (
);

FILL FILL_0__12835_ (
);

FILL FILL357200x19760 (
);

NAND2X1 _12700_ (
    .A(\datapath_1.alu_1.ALUInA [23]),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2265_)
);

OR2X2 _15592_ (
    .A(_4544_),
    .B(_4537_),
    .Y(_4545_)
);

AND2X2 _15172_ (
    .A(_4129_),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .Y(_4130_)
);

OR2X2 _9907_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_794__bF$buf0),
    .Y(_750_)
);

FILL FILL471200x247000 (
);

FILL FILL175560x128440 (
);

AND2X2 _13905_ (
    .A(_3336_),
    .B(_3335_),
    .Y(\datapath_1.alu_1.ALUInA [29])
);

AND2X2 _16797_ (
    .A(_4228__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_5731_)
);

OR2X2 _16377_ (
    .A(_5317_),
    .B(_5286_),
    .Y(_5318_)
);

FILL FILL_1__18460_ (
);

OR2X2 _11092_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_1388__bF$buf4),
    .Y(_1360_)
);

FILL FILL187720x69160 (
);

FILL FILL_0__17453_ (
);

FILL FILL_0__17033_ (
);

FILL FILL296400x167960 (
);

FILL FILL383800x172900 (
);

FILL FILL164160x69160 (
);

OR2X2 _9660_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_625_)
);

OR2X2 _9240_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_405_)
);

DFFSR _12297_ (
    .CLK(clk_bF$buf10),
    .D(_1917_[3]),
    .Q(\datapath_1.regfile_1.regOut[30] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL_1__14380_ (
);

FILL FILL_0__18658_ (
);

AND2X2 _18943_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_7845_)
);

AND2X2 _18523_ (
    .A(_6229__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_7431_)
);

AND2X2 _18103_ (
    .A(_6238__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_7018_)
);

FILL FILL_0__13793_ (
);

FILL FILL_0__13373_ (
);

FILL FILL397480x360620 (
);

FILL FILL290320x242060 (
);

FILL FILL_0__9700_ (
);

FILL FILL_1__15165_ (
);

AND2X2 _19308_ (
    .A(_6221__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_8204_)
);

DFFSR _14863_ (
    .CLK(clk_bF$buf98),
    .D(_3870_[11]),
    .Q(_2_[11]),
    .R(rst_bF$buf87),
    .S(vdd)
);

FILL FILL_0__14578_ (
);

FILL FILL_0__14158_ (
);

AND2X2 _14443_ (
    .A(_3721_),
    .B(_3720_),
    .Y(_3672_[24])
);

AND2X2 _14023_ (
    .A(_3344__bF$buf0),
    .B(gnd),
    .Y(_3439_)
);

FILL FILL_1__11085_ (
);

OR2X2 _15648_ (
    .A(_4599_),
    .B(_4596_),
    .Y(_4600_)
);

AND2X2 _15228_ (
    .A(_4133_),
    .B(_4171_),
    .Y(_4186_)
);

OR2X2 _10783_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_1256__bF$buf1),
    .Y(_1194_)
);

DFFSR _10363_ (
    .CLK(clk_bF$buf51),
    .D(_927_[4]),
    .Q(\datapath_1.regfile_1.regOut[15] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL_0__10078_ (
);

FILL FILL_0__16724_ (
);

FILL FILL_0__16304_ (
);

OR2X2 _19481_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_8356_)
);

AND2X2 _19061_ (
    .A(_6250__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_7961_)
);

FILL FILL385320x0 (
);

FILL FILL102600x340860 (
);

OR2X2 _8931_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_259_)
);

OR2X2 _8511_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_39_)
);

FILL FILL440040x14820 (
);

OR2X2 _11988_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_1817_)
);

OR2X2 _11568_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_1597_)
);

DFFSR _11148_ (
    .CLK(clk_bF$buf54),
    .D(_1323_[15]),
    .Q(\datapath_1.regfile_1.regOut[21] [15]),
    .R(rst_bF$buf24),
    .S(vdd)
);

FILL FILL_0__17929_ (
);

FILL FILL_0__17509_ (
);

FILL FILL_0__12644_ (
);

DFFSR _9716_ (
    .CLK(clk_bF$buf111),
    .D(_597_[2]),
    .Q(\datapath_1.regfile_1.regOut[10] [2]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL_1__8673_ (
);

FILL FILL_1__14016_ (
);

FILL FILL_0__13849_ (
);

AND2X2 _13714_ (
    .A(_3089__bF$buf0),
    .B(gnd),
    .Y(_3192_)
);

FILL FILL_0__13009_ (
);

AND2X2 _16186_ (
    .A(_5129_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd2 [14])
);

FILL FILL_1__9038_ (
);

FILL FILL_0__17682_ (
);

FILL FILL_0__17262_ (
);

FILL FILL_1__10356_ (
);

OR2X2 _14919_ (
    .A(\datapath_1.mux_pcsrc.dout [11]),
    .B(_4001__bF$buf4),
    .Y(_3959_)
);

FILL FILL254600x256880 (
);

FILL FILL_1__19474_ (
);

FILL FILL_0__10710_ (
);

AND2X2 _18752_ (
    .A(_6244__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_7657_)
);

AND2X2 _18332_ (
    .A(_6300__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_7243_)
);

FILL FILL_0__18047_ (
);

FILL FILL100320x202540 (
);

OR2X2 _10839_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_1231_)
);

OR2X2 _10419_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_1011_)
);

FILL FILL_1__15394_ (
);

DFFSR _19537_ (
    .CLK(clk_bF$buf98),
    .D(_8320_[14]),
    .Q(\datapath_1.regfile_1.regOut[0] [14]),
    .R(rst_bF$buf87),
    .S(vdd)
);

AND2X2 _19117_ (
    .A(_6247__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_8016_)
);

OR2X2 _14672_ (
    .A(vdd),
    .B(\datapath_1.a [15]),
    .Y(_3834_)
);

FILL FILL_0__14387_ (
);

OR2X2 _14252_ (
    .A(vdd),
    .B(ALUOut[4]),
    .Y(_3614_)
);

FILL FILL_1__13707_ (
);

FILL FILL430920x242060 (
);

FILL FILL448400x88920 (
);

FILL FILL500080x143260 (
);

AND2X2 _15877_ (
    .A(_4234__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_4825_)
);

AND2X2 _15457_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_4412_)
);

AND2X2 _15037_ (
    .A(_4025_),
    .B(_4022_),
    .Y(_4026_)
);

AND2X2 _10592_ (
    .A(_1106_),
    .B(_1105_),
    .Y(_1059_[23])
);

AND2X2 _10172_ (
    .A(_886_),
    .B(_885_),
    .Y(_861_[12])
);

FILL FILL_1__8729_ (
);

FILL FILL_0__16953_ (
);

FILL FILL_0__16533_ (
);

FILL FILL_0__16113_ (
);

FILL FILL261440x143260 (
);

FILL FILL407360x59280 (
);

OR2X2 _19290_ (
    .A(_8183_),
    .B(_8186_),
    .Y(_8187_)
);

FILL FILL298680x266760 (
);

OR2X2 _8740_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .B(_200__bF$buf1),
    .Y(_152_)
);

DFFSR _11797_ (
    .CLK(clk_bF$buf4),
    .D(_1653_[19]),
    .Q(\datapath_1.regfile_1.regOut[26] [19]),
    .R(rst_bF$buf20),
    .S(vdd)
);

FILL FILL_1__18325_ (
);

OR2X2 _11377_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_1520__bF$buf2),
    .Y(_1510_)
);

OR2X2 _17603_ (
    .A(_6493_),
    .B(_6525_),
    .Y(_6526_)
);

FILL FILL13680x321100 (
);

FILL FILL233320x276640 (
);

OR2X2 _9945_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_775_)
);

OR2X2 _9525_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_555_)
);

OR2X2 _9105_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_335_)
);

FILL FILL256120x360620 (
);

FILL FILL_1__14665_ (
);

AND2X2 _18808_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_7712_)
);

FILL FILL_0_BUFX2_insert251 (
);

FILL FILL_0_BUFX2_insert253 (
);

AND2X2 _13943_ (
    .A(_3352__bF$buf4),
    .B(\aluControl_1.inst [1]),
    .Y(_3371_)
);

FILL FILL_0__13658_ (
);

FILL FILL_0_BUFX2_insert254 (
);

FILL FILL_0__13238_ (
);

FILL FILL_0_BUFX2_insert255 (
);

OR2X2 _13523_ (
    .A(ALUOut[11]),
    .B(_3079__bF$buf3),
    .Y(_3037_)
);

AOI21X1 _13103_ (
    .A(_2271_),
    .B(_2272_),
    .C(_2501_),
    .Y(_2657_)
);

FILL FILL_0_BUFX2_insert256 (
);

FILL FILL_0_BUFX2_insert257 (
);

FILL FILL83600x207480 (
);

FILL FILL_0_BUFX2_insert258 (
);

FILL FILL438520x271700 (
);

FILL FILL368600x276640 (
);

FILL FILL_1__10165_ (
);

DFFSR _14728_ (
    .CLK(clk_bF$buf15),
    .D(_3804_[5]),
    .Q(\datapath_1.a [5]),
    .R(rst_bF$buf53),
    .S(vdd)
);

AND2X2 _14308_ (
    .A(_3651_),
    .B(_3650_),
    .Y(_3606_[22])
);

BUFX2 BUFX2_insert990 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf0)
);

BUFX2 BUFX2_insert991 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf4 )
);

BUFX2 BUFX2_insert992 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf3 )
);

BUFX2 BUFX2_insert993 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf2 )
);

BUFX2 BUFX2_insert994 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf1 )
);

BUFX2 BUFX2_insert995 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf0 )
);

BUFX2 BUFX2_insert996 (
    .A(_2157_),
    .Y(_2157__bF$buf3)
);

BUFX2 BUFX2_insert997 (
    .A(_2157_),
    .Y(_2157__bF$buf2)
);

BUFX2 BUFX2_insert998 (
    .A(_2157_),
    .Y(_2157__bF$buf1)
);

FILL FILL_0__15804_ (
);

BUFX2 BUFX2_insert999 (
    .A(_2157_),
    .Y(_2157__bF$buf0)
);

FILL FILL455240x187720 (
);

FILL FILL_0__18696_ (
);

AND2X2 _18981_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_7882_)
);

OR2X2 _18561_ (
    .A(_7461_),
    .B(_7468_),
    .Y(_7469_)
);

FILL FILL_0__18276_ (
);

AND2X2 _18141_ (
    .A(_6238__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_7055_)
);

FILL FILL_0__8797_ (
);

DFFSR _10648_ (
    .CLK(clk_bF$buf100),
    .D(_1059_[31]),
    .Q(\datapath_1.regfile_1.regOut[17] [31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL469680x148200 (
);

OR2X2 _10228_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .B(_926__bF$buf4),
    .Y(_924_)
);

FILL FILL_1__12731_ (
);

FILL FILL167200x4940 (
);

FILL FILL_0__11304_ (
);

AND2X2 _19346_ (
    .A(_6293__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_8242_)
);

DFFSR _14481_ (
    .CLK(clk_bF$buf78),
    .D(_3672_[16]),
    .Q(\datapath_1.Data [16]),
    .R(rst_bF$buf85),
    .S(vdd)
);

AND2X2 _14061_ (
    .A(_3350__bF$buf4),
    .B(_2_[20]),
    .Y(_3472_)
);

FILL FILL212040x296400 (
);

FILL FILL26600x148200 (
);

FILL FILL349600x222300 (
);

FILL FILL_0__12929_ (
);

FILL FILL_0__12509_ (
);

FILL FILL362520x217360 (
);

FILL FILL504640x251940 (
);

AND2X2 _15686_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_4637_)
);

AND2X2 _15266_ (
    .A(_4223__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_4224_)
);

FILL FILL_0__16762_ (
);

FILL FILL148200x335920 (
);

FILL FILL504640x0 (
);

FILL FILL_1__18974_ (
);

FILL FILL_1__18554_ (
);

AND2X2 _11186_ (
    .A(_1402_),
    .B(_1401_),
    .Y(_1389_[6])
);

FILL FILL_0__17547_ (
);

AND2X2 _17832_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_6751_)
);

AND2X2 _17412_ (
    .A(_6323__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_6337_)
);

FILL FILL_0__17127_ (
);

FILL FILL79800x330980 (
);

FILL FILL_0__12682_ (
);

FILL FILL_0__12262_ (
);

OR2X2 _9754_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_728__bF$buf1),
    .Y(_668_)
);

DFFSR _9334_ (
    .CLK(clk_bF$buf68),
    .D(_399_[7]),
    .Q(\datapath_1.regfile_1.regOut[7] [7]),
    .R(rst_bF$buf107),
    .S(vdd)
);

FILL FILL_1__14054_ (
);

OR2X2 _18617_ (
    .A(_7523_),
    .B(_7522_),
    .Y(_7524_)
);

FILL FILL_0__13887_ (
);

AND2X2 _13752_ (
    .A(_3081__bF$buf0),
    .B(ALUOut[23]),
    .Y(_3224_)
);

AND2X2 _13332_ (
    .A(_2872_),
    .B(_2408_),
    .Y(_2873_)
);

FILL FILL31920x158080 (
);

FILL FILL_1__15679_ (
);

FILL FILL_1__15259_ (
);

OR2X2 _14957_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [24]),
    .Y(_3984_)
);

FILL FILL115520x14820 (
);

OR2X2 _14537_ (
    .A(IRWrite_bF$buf4),
    .B(\datapath_1.PCJump [15]),
    .Y(_3764_)
);

AND2X2 _14117_ (
    .A(_3350__bF$buf2),
    .B(_2_[28]),
    .Y(_3520_)
);

FILL FILL229520x83980 (
);

OR2X2 _18790_ (
    .A(_7693_),
    .B(_7686_),
    .Y(_7694_)
);

FILL FILL227240x261820 (
);

FILL FILL_0__18085_ (
);

AND2X2 _18370_ (
    .A(_6229__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_7281_)
);

FILL FILL240160x256880 (
);

FILL FILL_1__11179_ (
);

FILL FILL364040x321100 (
);

DFFSR _10877_ (
    .CLK(clk_bF$buf90),
    .D(_1191_[2]),
    .Q(\datapath_1.regfile_1.regOut[19] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

AND2X2 _10457_ (
    .A(_1036_),
    .B(_1035_),
    .Y(_993_[21])
);

AND2X2 _10037_ (
    .A(_816_),
    .B(_815_),
    .Y(_795_[10])
);

FILL FILL_1__12960_ (
);

FILL FILL_1__12540_ (
);

FILL FILL_0__16818_ (
);

FILL FILL_0__11953_ (
);

AND2X2 _19155_ (
    .A(_6300__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_8054_)
);

AND2X2 _14290_ (
    .A(_3639_),
    .B(_3638_),
    .Y(_3606_[16])
);

OR2X2 _8605_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .B(_134__bF$buf3),
    .Y(_82_)
);

FILL FILL414200x54340 (
);

FILL FILL_0__12738_ (
);

INVX1 _12603_ (
    .A(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2168_)
);

FILL FILL435480x93860 (
);

OR2X2 _15495_ (
    .A(_4448_),
    .B(_4447_),
    .Y(_4449_)
);

OR2X2 _15075_ (
    .A(_4043_),
    .B(_4061_),
    .Y(_4062_)
);

FILL FILL115520x128440 (
);

FILL FILL_0__16151_ (
);

FILL FILL398240x340860 (
);

AND2X2 _13808_ (
    .A(_3081__bF$buf0),
    .B(ALUOut[31]),
    .Y(_3272_)
);

FILL FILL_0__17776_ (
);

AND2X2 _17641_ (
    .A(_6317__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_6563_)
);

AND2X2 _17221_ (
    .A(_4142__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_6148_)
);

FILL FILL_0__12491_ (
);

FILL FILL_0__12071_ (
);

DFFSR _9983_ (
    .CLK(clk_bF$buf45),
    .D(_729_[11]),
    .Q(\datapath_1.regfile_1.regOut[12] [11]),
    .R(rst_bF$buf57),
    .S(vdd)
);

AND2X2 _9563_ (
    .A(_580_),
    .B(_579_),
    .Y(_531_[24])
);

AND2X2 _9143_ (
    .A(_360_),
    .B(_359_),
    .Y(_333_[13])
);

FILL FILL_1__14283_ (
);

OR2X2 _18846_ (
    .A(_7748_),
    .B(_7747_),
    .Y(_7749_)
);

AND2X2 _18426_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_7336_)
);

FILL FILL_0_BUFX2_insert631 (
);

FILL FILL356440x202540 (
);

AND2X2 _18006_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_6922_)
);

FILL FILL_0_BUFX2_insert633 (
);

FILL FILL136040x286520 (
);

AND2X2 _13981_ (
    .A(_3344__bF$buf0),
    .B(gnd),
    .Y(_3403_)
);

FILL FILL_0_BUFX2_insert634 (
);

FILL FILL_0_BUFX2_insert635 (
);

FILL FILL_0__13276_ (
);

OR2X2 _13561_ (
    .A(IorD_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [24]),
    .Y(_3062_)
);

FILL FILL177840x14820 (
);

XOR2X1 _13141_ (
    .A(_2277_),
    .B(_2679_),
    .Y(_2693_)
);

FILL FILL_0_BUFX2_insert636 (
);

FILL FILL_0_BUFX2_insert637 (
);

FILL FILL_0_BUFX2_insert639 (
);

FILL FILL373920x212420 (
);

FILL FILL475760x83980 (
);

FILL FILL468160x158080 (
);

OR2X2 _14766_ (
    .A(\datapath_1.rd2 [3]),
    .B(_3935__bF$buf3),
    .Y(_3877_)
);

DFFSR _14346_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[10]),
    .Q(ALUOut[10]),
    .R(rst_bF$buf29),
    .S(vdd)
);

FILL FILL50160x365560 (
);

FILL FILL_0__15842_ (
);

FILL FILL_0__15422_ (
);

FILL FILL371640x286520 (
);

OR2X2 _10686_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_1149_)
);

OR2X2 _10266_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_929_)
);

FILL FILL_0__16627_ (
);

OR2X2 _16912_ (
    .A(_5840_),
    .B(_5843_),
    .Y(_5844_)
);

FILL FILL_0__11762_ (
);

FILL FILL_0__11342_ (
);

OR2X2 _19384_ (
    .A(_8278_),
    .B(_8277_),
    .Y(_8279_)
);

FILL FILL_0__19099_ (
);

DFFSR _8834_ (
    .CLK(clk_bF$buf25),
    .D(_135_[23]),
    .Q(\datapath_1.regfile_1.regOut[3] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL25840x143260 (
);

BUFX2 _8414_ (
    .A(_1_[22]),
    .Y(memoryAddress[22])
);

FILL FILL_1__18839_ (
);

FILL FILL_1__18419_ (
);

FILL FILL_1__13134_ (
);

FILL FILL504640x321100 (
);

FILL FILL248520x311220 (
);

FILL FILL_0__12967_ (
);

OR2X2 _12832_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2397_)
);

FILL FILL_0__12547_ (
);

OR2X2 _12412_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .B(_2048__bF$buf3),
    .Y(_2040_)
);

FILL FILL_0__12127_ (
);

FILL FILL329080x281580 (
);

OR2X2 _9619_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(_662__bF$buf3),
    .Y(_598_)
);

FILL FILL_0__16380_ (
);

OR2X2 _13617_ (
    .A(_3108_),
    .B(_3107_),
    .Y(_3109_)
);

FILL FILL_1__15700_ (
);

OR2X2 _16089_ (
    .A(_5018_),
    .B(_5033_),
    .Y(_5034_)
);

AND2X2 _17870_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_6788_)
);

AND2X2 _17450_ (
    .A(_6221__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_6375_)
);

FILL FILL_0__17165_ (
);

AND2X2 _17030_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_5960_)
);

OR2X2 _9792_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_693_)
);

OR2X2 _9372_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_473_)
);

FILL FILL_1__11620_ (
);

OR2X2 _18655_ (
    .A(_7559_),
    .B(_7560_),
    .Y(_7561_)
);

OR2X2 _18235_ (
    .A(_7140_),
    .B(_7147_),
    .Y(_7148_)
);

FILL FILL245480x4940 (
);

AND2X2 _13790_ (
    .A(_3087__bF$buf1),
    .B(\datapath_1.ALUResult [28]),
    .Y(_3257_)
);

FILL FILL_0__13085_ (
);

OR2X2 _13370_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2908_)
);

FILL FILL_0__19311_ (
);

FILL FILL386840x251940 (
);

FILL FILL_1__12825_ (
);

FILL FILL122360x108680 (
);

FILL FILL243200x281580 (
);

FILL FILL8360x261820 (
);

FILL FILL_0__9832_ (
);

FILL FILL_0__11818_ (
);

FILL FILL_0__9412_ (
);

DFFSR _14995_ (
    .CLK(clk_bF$buf62),
    .D(_3936_[14]),
    .Q(\datapath_1.mux_iord.din0 [14]),
    .R(rst_bF$buf18),
    .S(vdd)
);

AND2X2 _14575_ (
    .A(_3789_),
    .B(_3788_),
    .Y(_3738_[25])
);

OR2X2 _14155_ (
    .A(MemToReg_bF$buf1),
    .B(ALUOut[4]),
    .Y(_3548_)
);

FILL FILL278160x0 (
);

FILL FILL_0__15651_ (
);

FILL FILL_0__15231_ (
);

FILL FILL_1__17443_ (
);

DFFSR _10495_ (
    .CLK(clk_bF$buf48),
    .D(_993_[7]),
    .Q(\datapath_1.regfile_1.regOut[16] [7]),
    .R(rst_bF$buf14),
    .S(vdd)
);

OR2X2 _10075_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .B(_860__bF$buf1),
    .Y(_842_)
);

FILL FILL_1__17023_ (
);

AND2X2 _16721_ (
    .A(_4181__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_5656_)
);

FILL FILL_0__16016_ (
);

AND2X2 _16301_ (
    .A(_4241__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_5243_)
);

FILL FILL_0__11991_ (
);

FILL FILL_0__11571_ (
);

OR2X2 _19193_ (
    .A(_8083_),
    .B(_8090_),
    .Y(_8091_)
);

OR2X2 _8643_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_107_)
);

FILL FILL44840x123500 (
);

FILL FILL_1__13783_ (
);

OR2X2 _17926_ (
    .A(_6843_),
    .B(_6836_),
    .Y(_6844_)
);

AND2X2 _17506_ (
    .A(_6282__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_6430_)
);

FILL FILL_0__12776_ (
);

INVX1 _12641_ (
    .A(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2206_)
);

FILL FILL_0__12356_ (
);

AND2X2 _12221_ (
    .A(_1932_),
    .B(_1931_),
    .Y(_1917_[7])
);

FILL FILL361760x350740 (
);

DFFSR _9848_ (
    .CLK(clk_bF$buf36),
    .D(_663_[5]),
    .Q(\datapath_1.regfile_1.regOut[11] [5]),
    .R(rst_bF$buf78),
    .S(vdd)
);

AND2X2 _9428_ (
    .A(_510_),
    .B(_509_),
    .Y(_465_[22])
);

FILL FILL278920x360620 (
);

AND2X2 _9008_ (
    .A(_290_),
    .B(_289_),
    .Y(_267_[11])
);

FILL FILL16720x29640 (
);

FILL FILL417240x19760 (
);

FILL FILL_1__14148_ (
);

OR2X2 _13846_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [10]),
    .Y(_3297_)
);

OR2X2 _13426_ (
    .A(_2855_),
    .B(_2960_),
    .Y(_2961_)
);

OAI21X1 _13006_ (
    .A(_2321_),
    .B(_2503_),
    .C(_2565_),
    .Y(_2566_)
);

FILL FILL_0__14502_ (
);

FILL FILL_0__17394_ (
);

FILL FILL265240x98800 (
);

OR2X2 _9181_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .B(_398__bF$buf3),
    .Y(_386_)
);

FILL FILL149720x217360 (
);

FILL FILL_0__15707_ (
);

FILL FILL_0__10842_ (
);

OR2X2 _18884_ (
    .A(_7783_),
    .B(_7786_),
    .Y(_7787_)
);

FILL FILL_0__18599_ (
);

OR2X2 _18464_ (
    .A(_7372_),
    .B(_7369_),
    .Y(_7373_)
);

OR2X2 _18044_ (
    .A(_6959_),
    .B(_6958_),
    .Y(_6960_)
);

FILL FILL236360x128440 (
);

FILL FILL_1__17919_ (
);

FILL FILL272840x301340 (
);

FILL FILL_0__9641_ (
);

FILL FILL_0__11627_ (
);

DFFSR _11912_ (
    .CLK(clk_bF$buf70),
    .D(_1719_[5]),
    .Q(\datapath_1.regfile_1.regOut[27] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL_0__11207_ (
);

OR2X2 _19249_ (
    .A(_8144_),
    .B(_8145_),
    .Y(_8146_)
);

FILL FILL_0__14099_ (
);

OR2X2 _14384_ (
    .A(vdd),
    .B(\datapath_1.Data [5]),
    .Y(_3682_)
);

FILL FILL_0__15880_ (
);

FILL FILL_0__15040_ (
);

FILL FILL246240x9880 (
);

FILL FILL411920x39520 (
);

FILL FILL268280x19760 (
);

AND2X2 _15589_ (
    .A(_4130__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_4542_)
);

AND2X2 _15169_ (
    .A(_4126_),
    .B(\datapath_1.PCJump [18]),
    .Y(_4127_)
);

FILL FILL331360x345800 (
);

FILL FILL_1__17672_ (
);

FILL FILL_0__16665_ (
);

OR2X2 _16950_ (
    .A(_5878_),
    .B(_5881_),
    .Y(_5882_)
);

AND2X2 _16530_ (
    .A(_4167__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_5468_)
);

FILL FILL_0__16245_ (
);

OR2X2 _16110_ (
    .A(_5053_),
    .B(_5054_),
    .Y(_5055_)
);

FILL FILL_0__11380_ (
);

OR2X2 _8872_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .B(_266__bF$buf0),
    .Y(_220_)
);

BUFX2 _8452_ (
    .A(_2_[28]),
    .Y(memoryWriteData[28])
);

FILL FILL231800x192660 (
);

OR2X2 _11089_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_1388__bF$buf1),
    .Y(_1358_)
);

FILL FILL_1__13172_ (
);

AND2X2 _17735_ (
    .A(_6655_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd1 [5])
);

OR2X2 _17315_ (
    .A(_6234_),
    .B(_6240_),
    .Y(_6241_)
);

NAND2X1 _12870_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2435_)
);

FILL FILL423320x281580 (
);

DFFSR _12450_ (
    .CLK(clk_bF$buf14),
    .D(_1983_[27]),
    .Q(\datapath_1.regfile_1.regOut[31] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

OR2X2 _12030_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_1845_)
);

FILL FILL_0__18811_ (
);

OR2X2 _9657_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_623_)
);

OR2X2 _9237_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_403_)
);

FILL FILL323000x375440 (
);

FILL FILL114760x261820 (
);

FILL FILL_0__8912_ (
);

FILL FILL145920x247000 (
);

FILL FILL215080x148200 (
);

AND2X2 _13655_ (
    .A(_3084__bF$buf1),
    .B(\datapath_1.PCJump [9]),
    .Y(_3141_)
);

OR2X2 _13235_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2781_)
);

FILL FILL267520x4940 (
);

FILL FILL_1__10297_ (
);

FILL FILL42560x83980 (
);

FILL FILL_1__16523_ (
);

FILL FILL51680x103740 (
);

FILL FILL418760x266760 (
);

OR2X2 _15801_ (
    .A(_4719_),
    .B(_4750_),
    .Y(_4751_)
);

FILL FILL_0__15516_ (
);

FILL FILL32680x261820 (
);

AND2X2 _18693_ (
    .A(_6238__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_7599_)
);

AND2X2 _18273_ (
    .A(_6328__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_7185_)
);

FILL FILL299440x316160 (
);

FILL FILL_1__17308_ (
);

FILL FILL504640x88920 (
);

FILL FILL_0__9450_ (
);

OR2X2 _11721_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_1679_)
);

FILL FILL_0__11436_ (
);

FILL FILL_0__9030_ (
);

OR2X2 _11301_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_1459_)
);

OR2X2 _19478_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_8354_)
);

AND2X2 _19058_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_7958_)
);

AND2X2 _14193_ (
    .A(_3573_),
    .B(_3572_),
    .Y(\datapath_1.mux_wd3.dout [16])
);

OR2X2 _8928_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_257_)
);

OR2X2 _8508_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_37_)
);

FILL FILL_1__13648_ (
);

AND2X2 _12926_ (
    .A(_2490_),
    .B(_2163_),
    .Y(_2491_)
);

NOR2X1 _12506_ (
    .A(_2101_),
    .B(_2102_),
    .Y(RegDst)
);

FILL FILL315400x256880 (
);

FILL FILL_1_BUFX2_insert566 (
);

FILL FILL_1_BUFX2_insert568 (
);

OR2X2 _15398_ (
    .A(_4352_),
    .B(_4353_),
    .Y(_4354_)
);

FILL FILL480320x34580 (
);

FILL FILL370880x54340 (
);

FILL FILL_1__17061_ (
);

FILL FILL_0__16894_ (
);

FILL FILL_0__16474_ (
);

AND2X2 _8681_ (
    .A(_132_),
    .B(_131_),
    .Y(_69_[31])
);

FILL FILL253840x93860 (
);

FILL FILL183160x69160 (
);

BUFX2 BUFX2_insert230 (
    .A(_4187_),
    .Y(_4187__bF$buf3)
);

BUFX2 BUFX2_insert231 (
    .A(_4187_),
    .Y(_4187__bF$buf2)
);

BUFX2 BUFX2_insert232 (
    .A(_4187_),
    .Y(_4187__bF$buf1)
);

BUFX2 BUFX2_insert233 (
    .A(_4187_),
    .Y(_4187__bF$buf0)
);

BUFX2 BUFX2_insert234 (
    .A(_1982_),
    .Y(_1982__bF$buf4)
);

AND2X2 _17964_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_6881_)
);

FILL FILL_0__17679_ (
);

AND2X2 _17544_ (
    .A(_6287__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_6467_)
);

FILL FILL_0__17259_ (
);

BUFX2 BUFX2_insert235 (
    .A(_1982_),
    .Y(_1982__bF$buf3)
);

BUFX2 BUFX2_insert236 (
    .A(_1982_),
    .Y(_1982__bF$buf2)
);

AND2X2 _17124_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_6053_)
);

BUFX2 BUFX2_insert237 (
    .A(_1982_),
    .Y(_1982__bF$buf1)
);

BUFX2 BUFX2_insert238 (
    .A(_1982_),
    .Y(_1982__bF$buf0)
);

FILL FILL_0__12394_ (
);

BUFX2 BUFX2_insert239 (
    .A(_6236_),
    .Y(_6236__bF$buf4)
);

FILL FILL177840x128440 (
);

OR2X2 _9886_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .B(_794__bF$buf4),
    .Y(_736_)
);

DFFSR _9466_ (
    .CLK(clk_bF$buf30),
    .D(_465_[10]),
    .Q(\datapath_1.regfile_1.regOut[8] [10]),
    .R(rst_bF$buf64),
    .S(vdd)
);

OR2X2 _9046_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .B(_332__bF$buf0),
    .Y(_316_)
);

FILL FILL283480x202540 (
);

FILL FILL484120x34580 (
);

FILL FILL158840x286520 (
);

FILL FILL_0__8721_ (
);

FILL FILL7600x54340 (
);

AND2X2 _18749_ (
    .A(_6312__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_7654_)
);

AND2X2 _18329_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_7240_)
);

AND2X2 _13884_ (
    .A(_3322_),
    .B(_3321_),
    .Y(\datapath_1.alu_1.ALUInA [22])
);

FILL FILL_0__13599_ (
);

AND2X2 _13464_ (
    .A(_2996_),
    .B(_2878_),
    .Y(_2997_)
);

FILL FILL_0__13179_ (
);

AND2X2 _13044_ (
    .A(_2600_),
    .B(_2302_),
    .Y(_2601_)
);

FILL FILL_0__19405_ (
);

FILL FILL_0__14540_ (
);

FILL FILL_0__14120_ (
);

FILL FILL281960x370500 (
);

FILL FILL408120x158080 (
);

FILL FILL163400x39520 (
);

FILL FILL_0__9926_ (
);

FILL FILL_0__9506_ (
);

FILL FILL505400x301340 (
);

OR2X2 _14669_ (
    .A(vdd),
    .B(\datapath_1.a [14]),
    .Y(_3832_)
);

OR2X2 _14249_ (
    .A(vdd),
    .B(ALUOut[3]),
    .Y(_3612_)
);

FILL FILL400520x123500 (
);

FILL FILL338200x49400 (
);

FILL FILL_0__15745_ (
);

AND2X2 _15610_ (
    .A(_4562_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd2 [5])
);

FILL FILL_0__10460_ (
);

FILL FILL_0__10040_ (
);

AND2X2 _18082_ (
    .A(_6229__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_6997_)
);

FILL FILL399760x360620 (
);

FILL FILL292600x242060 (
);

AND2X2 _10589_ (
    .A(_1104_),
    .B(_1103_),
    .Y(_1059_[22])
);

FILL FILL_1__17537_ (
);

AND2X2 _10169_ (
    .A(_884_),
    .B(_883_),
    .Y(_861_[11])
);

FILL FILL161120x350740 (
);

OR2X2 _16815_ (
    .A(_5745_),
    .B(_5748_),
    .Y(_5749_)
);

FILL FILL207480x256880 (
);

FILL FILL152760x227240 (
);

OR2X2 _11950_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_1850__bF$buf3),
    .Y(_1792_)
);

DFFSR _11530_ (
    .CLK(clk_bF$buf107),
    .D(_1521_[10]),
    .Q(\datapath_1.regfile_1.regOut[24] [10]),
    .R(rst_bF$buf95),
    .S(vdd)
);

OR2X2 _11110_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .B(_1388__bF$buf1),
    .Y(_1372_)
);

AND2X2 _19287_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_8184_)
);

FILL FILL167200x39520 (
);

OR2X2 _8737_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .B(_200__bF$buf3),
    .Y(_150_)
);

FILL FILL9120x158080 (
);

NAND2X1 _12735_ (
    .A(\datapath_1.alu_1.ALUInA [19]),
    .B(_2299_),
    .Y(_2300_)
);

DFFSR _12315_ (
    .CLK(clk_bF$buf43),
    .D(_1917_[21]),
    .Q(\datapath_1.regfile_1.regOut[30] [21]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL_0__13811_ (
);

FILL FILL9880x143260 (
);

FILL FILL_0__16283_ (
);

FILL FILL446120x64220 (
);

FILL FILL_1__9420_ (
);

OR2X2 _8490_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_25_)
);

FILL FILL130720x281580 (
);

FILL FILL_1__18495_ (
);

FILL FILL_0__17488_ (
);

OR2X2 _17773_ (
    .A(_6689_),
    .B(_6692_),
    .Y(_6693_)
);

FILL FILL_0__17068_ (
);

NAND3X1 _17353_ (
    .A(_6203_),
    .B(_6201_),
    .C(_6227_),
    .Y(_6279_)
);

FILL FILL486400x286520 (
);

AND2X2 _9695_ (
    .A(_648_),
    .B(_647_),
    .Y(_597_[25])
);

AND2X2 _9275_ (
    .A(_428_),
    .B(_427_),
    .Y(_399_[14])
);

FILL FILL_0__8530_ (
);

OR2X2 _10801_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_1256__bF$buf4),
    .Y(_1206_)
);

AND2X2 _18978_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_7879_)
);

AND2X2 _18558_ (
    .A(_6317__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_7466_)
);

OR2X2 _18138_ (
    .A(_7050_),
    .B(_7051_),
    .Y(_7052_)
);

AND2X2 _13693_ (
    .A(_3089__bF$buf1),
    .B(gnd),
    .Y(_3174_)
);

OR2X2 _13273_ (
    .A(_2387__bF$buf3),
    .B(_2816_),
    .Y(_2817_)
);

FILL FILL131480x247000 (
);

OR2X2 _14898_ (
    .A(\datapath_1.mux_pcsrc.dout [4]),
    .B(_4001__bF$buf4),
    .Y(_3945_)
);

DFFSR _14478_ (
    .CLK(clk_bF$buf23),
    .D(_3672_[13]),
    .Q(\datapath_1.Data [13]),
    .R(rst_bF$buf33),
    .S(vdd)
);

AND2X2 _14058_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3469_)
);

FILL FILL_1__16561_ (
);

FILL FILL_1__16141_ (
);

FILL FILL_0__15134_ (
);

FILL FILL205200x0 (
);

FILL FILL102600x202540 (
);

FILL FILL348840x0 (
);

OR2X2 _10398_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_997_)
);

FILL FILL_0__16759_ (
);

AND2X2 _16624_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_5561_)
);

FILL FILL_0__16339_ (
);

OR2X2 _16204_ (
    .A(_5145_),
    .B(_5146_),
    .Y(_5147_)
);

FILL FILL_0__11894_ (
);

FILL FILL266000x345800 (
);

OR2X2 _19096_ (
    .A(_7988_),
    .B(_7995_),
    .Y(_7996_)
);

FILL FILL_0__17700_ (
);

DFFSR _8966_ (
    .CLK(clk_bF$buf109),
    .D(_201_[26]),
    .Q(\datapath_1.regfile_1.regOut[4] [26]),
    .R(rst_bF$buf84),
    .S(vdd)
);

AND2X2 _8546_ (
    .A(_62_),
    .B(_61_),
    .Y(_3_[29])
);

FILL FILL_1__13266_ (
);

FILL FILL169480x187720 (
);

OR2X2 _17829_ (
    .A(_6747_),
    .B(_6740_),
    .Y(_6748_)
);

OR2X2 _17409_ (
    .A(_6269_),
    .B(_6334_),
    .Y(_6335_)
);

AND2X2 _12964_ (
    .A(_2526_),
    .B(_2520_),
    .Y(_2527_)
);

FILL FILL_0__12259_ (
);

OR2X2 _12544_ (
    .A(\control_1.op [2]),
    .B(\control_1.op [3]),
    .Y(_2133_)
);

OR2X2 _12124_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .B(_1916__bF$buf3),
    .Y(_1888_)
);

FILL FILL_1_BUFX2_insert946 (
);

FILL FILL_1_BUFX2_insert948 (
);

FILL FILL_0__18905_ (
);

FILL FILL_0__13620_ (
);

FILL FILL_0__13200_ (
);

FILL FILL_0__16092_ (
);

AND2X2 _13749_ (
    .A(_3089__bF$buf2),
    .B(gnd),
    .Y(_3222_)
);

NAND2X1 _13329_ (
    .A(_2869_),
    .B(_2867_),
    .Y(_2870_)
);

FILL FILL_0__14825_ (
);

FILL FILL_0__14405_ (
);

FILL FILL15960x321100 (
);

BUFX2 BUFX2_insert610 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf29)
);

BUFX2 BUFX2_insert611 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf28)
);

BUFX2 BUFX2_insert612 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf27)
);

BUFX2 BUFX2_insert613 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf26)
);

BUFX2 BUFX2_insert614 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf25)
);

AND2X2 _17582_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_6505_)
);

BUFX2 BUFX2_insert615 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf24)
);

BUFX2 BUFX2_insert616 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf23)
);

AND2X2 _17162_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_6090_)
);

BUFX2 BUFX2_insert617 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf22)
);

BUFX2 BUFX2_insert618 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf21)
);

BUFX2 BUFX2_insert619 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf20)
);

FILL FILL303240x44460 (
);

FILL FILL258400x360620 (
);

DFFSR _9084_ (
    .CLK(clk_bF$buf112),
    .D(_267_[15]),
    .Q(\datapath_1.regfile_1.regOut[5] [15]),
    .R(rst_bF$buf113),
    .S(vdd)
);

FILL FILL_1__11752_ (
);

FILL FILL213560x79040 (
);

FILL FILL_0__10325_ (
);

AND2X2 _10610_ (
    .A(_1118_),
    .B(_1117_),
    .Y(_1059_[29])
);

AND2X2 _18787_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_7691_)
);

AND2X2 _18367_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_7278_)
);

AND2X2 _13082_ (
    .A(_2636_),
    .B(_2270_),
    .Y(_2637_)
);

FILL FILL_0__19443_ (
);

FILL FILL_0__19023_ (
);

FILL FILL212800x301340 (
);

FILL FILL_1__12117_ (
);

FILL FILL_0__9964_ (
);

FILL FILL_0__9544_ (
);

OR2X2 _11815_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_1784__bF$buf3),
    .Y(_1722_)
);

FILL FILL237880x14820 (
);

FILL FILL212040x207480 (
);

AND2X2 _14287_ (
    .A(_3637_),
    .B(_3636_),
    .Y(_3606_[15])
);

FILL FILL_1__16790_ (
);

FILL FILL_0__15783_ (
);

FILL FILL_0__15363_ (
);

FILL FILL441560x29640 (
);

FILL FILL_1__8920_ (
);

FILL FILL242440x163020 (
);

FILL FILL217360x79040 (
);

FILL FILL234080x29640 (
);

FILL FILL207480x326040 (
);

FILL FILL159600x34580 (
);

FILL FILL_0__16988_ (
);

FILL FILL_0__16568_ (
);

AND2X2 _16853_ (
    .A(_4151__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_5786_)
);

AND2X2 _16433_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_5373_)
);

FILL FILL_0__16148_ (
);

AND2X2 _16013_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_4959_)
);

FILL FILL214320x296400 (
);

OR2X2 _8775_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_175_)
);

FILL FILL44840x39520 (
);

AND2X2 _17638_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_6560_)
);

AND2X2 _17218_ (
    .A(_4189__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_6145_)
);

OR2X2 _12773_ (
    .A(_2337_),
    .B(_2317_),
    .Y(_2338_)
);

FILL FILL_0__12488_ (
);

AND2X2 _12353_ (
    .A(_2000_),
    .B(_1999_),
    .Y(_1983_[8])
);

FILL FILL_0__12068_ (
);

FILL FILL_1__19301_ (
);

FILL FILL377720x163020 (
);

FILL FILL390640x158080 (
);

FILL FILL365560x44460 (
);

FILL FILL218880x88920 (
);

AND2X2 _13978_ (
    .A(_3352__bF$buf4),
    .B(\datapath_1.PCJump [8]),
    .Y(_3401_)
);

OR2X2 _13558_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [23]),
    .Y(_3060_)
);

INVX1 _13138_ (
    .A(_2676_),
    .Y(_2690_)
);

FILL FILL_1__15641_ (
);

FILL FILL117800x64220 (
);

FILL FILL_0__14634_ (
);

FILL FILL_0__14214_ (
);

AND2X2 _17391_ (
    .A(_6215_),
    .B(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_6317_)
);

FILL FILL_1__16006_ (
);

FILL FILL_0__15839_ (
);

OR2X2 _15704_ (
    .A(_4647_),
    .B(_4654_),
    .Y(_4655_)
);

FILL FILL194560x34580 (
);

FILL FILL_0__10974_ (
);

FILL FILL_0__10134_ (
);

AND2X2 _18596_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_7503_)
);

OR2X2 _18176_ (
    .A(_7088_),
    .B(_7089_),
    .Y(_7090_)
);

FILL FILL7600x345800 (
);

FILL FILL231040x321100 (
);

FILL FILL_0__19252_ (
);

FILL FILL225720x340860 (
);

FILL FILL_1__12766_ (
);

AND2X2 _16909_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_5841_)
);

FILL FILL_0__9773_ (
);

AND2X2 _11624_ (
    .A(_1634_),
    .B(_1633_),
    .Y(_1587_[23])
);

FILL FILL_0__11339_ (
);

FILL FILL411920x355680 (
);

AND2X2 _11204_ (
    .A(_1414_),
    .B(_1413_),
    .Y(_1389_[12])
);

FILL FILL408880x306280 (
);

AND2X2 _14096_ (
    .A(_3350__bF$buf4),
    .B(_2_[25]),
    .Y(_3502_)
);

FILL FILL_0__12700_ (
);

FILL FILL168720x291460 (
);

FILL FILL342000x29640 (
);

FILL FILL232560x49400 (
);

FILL FILL_0__15592_ (
);

OR2X2 _12829_ (
    .A(_2392_),
    .B(_2393_),
    .Y(_2394_)
);

FILL FILL366320x321100 (
);

OR2X2 _12409_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .B(_2048__bF$buf1),
    .Y(_2038_)
);

FILL FILL_1__14912_ (
);

FILL FILL_0__13905_ (
);

FILL FILL_0__16797_ (
);

OR2X2 _16662_ (
    .A(_5597_),
    .B(_5596_),
    .Y(_5598_)
);

OR2X2 _16242_ (
    .A(_5183_),
    .B(_5184_),
    .Y(_5185_)
);

FILL FILL_0__11092_ (
);

FILL FILL437000x54340 (
);

FILL FILL171000x19760 (
);

DFFSR _8584_ (
    .CLK(clk_bF$buf46),
    .D(_3_[31]),
    .Q(\datapath_1.regfile_1.regOut[1] [31]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL86640x291460 (
);

FILL FILL377720x256880 (
);

AND2X2 _17867_ (
    .A(_6250__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_6785_)
);

OR2X2 _17447_ (
    .A(_6370_),
    .B(_6371_),
    .Y(_6372_)
);

AND2X2 _17027_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_5957_)
);

OR2X2 _12582_ (
    .A(\control_1.next [3]),
    .B(_2145_),
    .Y(_2152_)
);

OR2X2 _12162_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_1913_)
);

FILL FILL_0__18943_ (
);

FILL FILL_0__18523_ (
);

FILL FILL_0__18103_ (
);

OR2X2 _9789_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_691_)
);

OR2X2 _9369_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_471_)
);

FILL FILL_0__8624_ (
);

FILL FILL_1__14089_ (
);

AND2X2 _13787_ (
    .A(_3081__bF$buf1),
    .B(ALUOut[28]),
    .Y(_3254_)
);

INVX1 _13367_ (
    .A(_2905_),
    .Y(\datapath_1.ALUResult [5])
);

FILL FILL_1__15030_ (
);

FILL FILL_0__19308_ (
);

FILL FILL287280x83980 (
);

FILL FILL166440x153140 (
);

FILL FILL_0__14023_ (
);

FILL FILL221920x370500 (
);

CLKBUF1 CLKBUF1_insert150 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf73)
);

CLKBUF1 CLKBUF1_insert151 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf72)
);

CLKBUF1 CLKBUF1_insert152 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf71)
);

CLKBUF1 CLKBUF1_insert153 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf70)
);

CLKBUF1 CLKBUF1_insert154 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert155 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf68)
);

CLKBUF1 CLKBUF1_insert156 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf67)
);

CLKBUF1 CLKBUF1_insert157 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert158 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf65)
);

CLKBUF1 CLKBUF1_insert159 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf64)
);

FILL FILL_1__16655_ (
);

FILL FILL_1__11370_ (
);

OR2X2 _15933_ (
    .A(_4879_),
    .B(_4878_),
    .Y(_4880_)
);

FILL FILL_0__15648_ (
);

OR2X2 _15513_ (
    .A(_4451_),
    .B(_4466_),
    .Y(_4467_)
);

FILL FILL_0__15228_ (
);

FILL FILL_0__10783_ (
);

FILL FILL_0__19481_ (
);

FILL FILL71440x207480 (
);

FILL FILL269800x365560 (
);

AND2X2 _16718_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_5653_)
);

FILL FILL_1__18801_ (
);

OR2X2 _11853_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_1747_)
);

FILL FILL_0__9162_ (
);

OR2X2 _11433_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_1527_)
);

DFFSR _11013_ (
    .CLK(clk_bF$buf113),
    .D(_1257_[9]),
    .Q(\datapath_1.regfile_1.regOut[20] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

FILL FILL430920x335920 (
);

FILL FILL133000x49400 (
);

FILL FILL115520x311220 (
);

FILL FILL373920x286520 (
);

FILL FILL56240x286520 (
);

FILL FILL443080x187720 (
);

FILL FILL301720x326040 (
);

INVX1 _12638_ (
    .A(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2203_)
);

AND2X2 _12218_ (
    .A(_1930_),
    .B(_1929_),
    .Y(_1917_[6])
);

FILL FILL38000x88920 (
);

FILL FILL_0__13714_ (
);

AND2X2 _16891_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_5823_)
);

FILL FILL_0__16186_ (
);

OR2X2 _16471_ (
    .A(_5409_),
    .B(_5406_),
    .Y(_5410_)
);

AND2X2 _16051_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_4997_)
);

FILL FILL386080x0 (
);

FILL FILL_1__9323_ (
);

FILL FILL10640x227240 (
);

FILL FILL_1__15506_ (
);

BUFX2 _8393_ (
    .A(_1_[1]),
    .Y(memoryAddress[1])
);

FILL FILL_0__14919_ (
);

FILL FILL87400x0 (
);

OR2X2 _17676_ (
    .A(_6596_),
    .B(_6595_),
    .Y(_6597_)
);

OR2X2 _17256_ (
    .A(_6182_),
    .B(_6175_),
    .Y(_6183_)
);

OR2X2 _12391_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .B(_2048__bF$buf3),
    .Y(_2026_)
);

FILL FILL_0__18752_ (
);

DFFSR _9598_ (
    .CLK(clk_bF$buf13),
    .D(_531_[13]),
    .Q(\datapath_1.regfile_1.regOut[9] [13]),
    .R(rst_bF$buf90),
    .S(vdd)
);

OR2X2 _9178_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .B(_398__bF$buf4),
    .Y(_384_)
);

FILL FILL_1__11426_ (
);

FILL FILL_0__8853_ (
);

OR2X2 _10704_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_1161_)
);

FILL FILL_0__10419_ (
);

FILL FILL_0_BUFX2_insert980 (
);

FILL FILL_0_BUFX2_insert982 (
);

FILL FILL373160x301340 (
);

FILL FILL_0_BUFX2_insert984 (
);

FILL FILL136040x335920 (
);

OR2X2 _13596_ (
    .A(_3090_),
    .B(_3088_),
    .Y(_3091_)
);

AND2X2 _13176_ (
    .A(_2725_),
    .B(_2723_),
    .Y(_2726_)
);

FILL FILL_0_BUFX2_insert986 (
);

FILL FILL_0_BUFX2_insert988 (
);

FILL FILL_0_BUFX2_insert989 (
);

AND2X2 _19402_ (
    .A(_6236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_8297_)
);

FILL FILL_0__19117_ (
);

FILL FILL_0__14252_ (
);

FILL FILL390640x311220 (
);

FILL FILL153520x345800 (
);

DFFSR _11909_ (
    .CLK(clk_bF$buf17),
    .D(_1719_[2]),
    .Q(\datapath_1.regfile_1.regOut[27] [2]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL_0__15877_ (
);

FILL FILL433200x98800 (
);

AND2X2 _15742_ (
    .A(_4210__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_4692_)
);

FILL FILL_0__15457_ (
);

AND2X2 _15322_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_4279_)
);

FILL FILL_0__10592_ (
);

FILL FILL415720x69160 (
);

FILL FILL_0__10172_ (
);

FILL FILL501600x291460 (
);

FILL FILL489440x138320 (
);

FILL FILL288800x345800 (
);

AND2X2 _16947_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_5879_)
);

OR2X2 _16527_ (
    .A(_5464_),
    .B(_5463_),
    .Y(_5465_)
);

OR2X2 _16107_ (
    .A(_5050_),
    .B(_5051_),
    .Y(_5052_)
);

FILL FILL_0__9391_ (
);

DFFSR _11662_ (
    .CLK(clk_bF$buf63),
    .D(_1587_[13]),
    .Q(\datapath_1.regfile_1.regOut[25] [13]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL_0__11377_ (
);

OR2X2 _11242_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .B(_1454__bF$buf2),
    .Y(_1440_)
);

OR2X2 _8869_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .B(_266__bF$buf2),
    .Y(_218_)
);

FILL FILL262200x88920 (
);

FILL FILL15960x14820 (
);

BUFX2 _8449_ (
    .A(_2_[25]),
    .Y(memoryWriteData[25])
);

OR2X2 _9810_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_705_)
);

FILL FILL_1__13589_ (
);

AOI22X1 _12867_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .C(\datapath_1.alu_1.ALUInB [8]),
    .D(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2432_)
);

DFFSR _12447_ (
    .CLK(clk_bF$buf6),
    .D(_1983_[24]),
    .Q(\datapath_1.regfile_1.regOut[31] [24]),
    .R(rst_bF$buf31),
    .S(vdd)
);

OR2X2 _12027_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_1843_)
);

FILL FILL145920x360620 (
);

FILL FILL_0__18808_ (
);

FILL FILL259920x108680 (
);

FILL FILL_0__13103_ (
);

FILL FILL456000x123500 (
);

OR2X2 _16280_ (
    .A(_5214_),
    .B(_5221_),
    .Y(_5222_)
);

FILL FILL95000x163020 (
);

FILL FILL_1__10450_ (
);

FILL FILL_0__14308_ (
);

OR2X2 _17485_ (
    .A(_6407_),
    .B(_6408_),
    .Y(_6409_)
);

AND2X2 _17065_ (
    .A(_4214__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_5995_)
);

FILL FILL_0__18561_ (
);

FILL FILL_0__18141_ (
);

FILL FILL_0__8662_ (
);

OR2X2 _10933_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .B(_1322__bF$buf2),
    .Y(_1274_)
);

FILL FILL_0__10228_ (
);

DFFSR _10513_ (
    .CLK(clk_bF$buf16),
    .D(_993_[25]),
    .Q(\datapath_1.regfile_1.regOut[16] [25]),
    .R(rst_bF$buf76),
    .S(vdd)
);

FILL FILL_0__19346_ (
);

AND2X2 _19211_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_8109_)
);

FILL FILL198360x172900 (
);

FILL FILL_0__14061_ (
);

FILL FILL_0__9447_ (
);

OR2X2 _11718_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_1677_)
);

FILL FILL107160x370500 (
);

FILL FILL120080x365560 (
);

FILL FILL498560x256880 (
);

FILL FILL321480x118560 (
);

OR2X2 _15971_ (
    .A(_4916_),
    .B(_4917_),
    .Y(_4918_)
);

FILL FILL_0__15686_ (
);

FILL FILL_0__15266_ (
);

AND2X2 _15551_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_4504_)
);

NOR2X1 _15131_ (
    .A(_4032_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.regfile_1.regEn [15])
);

FILL FILL344280x202540 (
);

FILL FILL_1__17478_ (
);

AND2X2 _16756_ (
    .A(_4241__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_5691_)
);

OR2X2 _16336_ (
    .A(_5273_),
    .B(_5276_),
    .Y(_5277_)
);

AND2X2 _11891_ (
    .A(_1772_),
    .B(_1771_),
    .Y(_1719_[26])
);

AND2X2 _11471_ (
    .A(_1552_),
    .B(_1551_),
    .Y(_1521_[15])
);

FILL FILL_0__11186_ (
);

AND2X2 _11051_ (
    .A(_1332_),
    .B(_1331_),
    .Y(_1323_[4])
);

FILL FILL283480x59280 (
);

FILL FILL351120x172900 (
);

FILL FILL_0__17412_ (
);

FILL FILL342760x370500 (
);

AND2X2 _8678_ (
    .A(_130_),
    .B(_129_),
    .Y(_69_[30])
);

FILL FILL291840x217360 (
);

FILL FILL434720x39520 (
);

AND2X2 _12676_ (
    .A(_2238_),
    .B(_2240_),
    .Y(_2241_)
);

OR2X2 _12256_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .B(_1982__bF$buf3),
    .Y(_1956_)
);

OR2X2 _18902_ (
    .A(_7788_),
    .B(_7804_),
    .Y(_7805_)
);

FILL FILL_0__18617_ (
);

FILL FILL259160x286520 (
);

FILL FILL_0__13752_ (
);

FILL FILL_0__13332_ (
);

FILL FILL216600x182780 (
);

FILL FILL354920x54340 (
);

FILL FILL_1__9781_ (
);

FILL FILL437000x4940 (
);

FILL FILL_1__15124_ (
);

FILL FILL_0__14957_ (
);

OR2X2 _14822_ (
    .A(vdd),
    .B(_2_[22]),
    .Y(_3914_)
);

FILL FILL_0__14537_ (
);

FILL FILL13680x143260 (
);

OR2X2 _14402_ (
    .A(vdd),
    .B(\datapath_1.Data [11]),
    .Y(_3694_)
);

FILL FILL421800x93860 (
);

AND2X2 _17294_ (
    .A(_6203_),
    .B(_6219_),
    .Y(_6220_)
);

FILL FILL405080x316160 (
);

FILL FILL_0__18790_ (
);

FILL FILL_0__18370_ (
);

FILL FILL_1__16329_ (
);

OR2X2 _15607_ (
    .A(_4559_),
    .B(_4552_),
    .Y(_4560_)
);

FILL FILL_0__8891_ (
);

FILL FILL_0__8471_ (
);

FILL FILL_0__10457_ (
);

AND2X2 _10742_ (
    .A(_1186_),
    .B(_1185_),
    .Y(_1125_[30])
);

AND2X2 _10322_ (
    .A(_966_),
    .B(_965_),
    .Y(_927_[19])
);

FILL FILL_0__10037_ (
);

FILL FILL203680x172900 (
);

OR2X2 _18499_ (
    .A(_7406_),
    .B(_7407_),
    .Y(_7408_)
);

AND2X2 _18079_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_6994_)
);

FILL FILL88920x83980 (
);

FILL FILL253080x227240 (
);

OR2X2 _19440_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8329_)
);

AND2X2 _19020_ (
    .A(_6315__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_7921_)
);

FILL FILL180120x59280 (
);

FILL FILL_0__14290_ (
);

FILL FILL_0__9676_ (
);

FILL FILL_0__9256_ (
);

OR2X2 _11947_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .B(_1850__bF$buf2),
    .Y(_1790_)
);

DFFSR _11527_ (
    .CLK(clk_bF$buf48),
    .D(_1521_[7]),
    .Q(\datapath_1.regfile_1.regOut[24] [7]),
    .R(rst_bF$buf21),
    .S(vdd)
);

OR2X2 _11107_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .B(_1388__bF$buf0),
    .Y(_1370_)
);

FILL FILL425600x93860 (
);

FILL FILL53960x103740 (
);

FILL FILL48640x237120 (
);

FILL FILL_0__12603_ (
);

FILL FILL_1__16082_ (
);

AND2X2 _15780_ (
    .A(_4225__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_4730_)
);

FILL FILL_0__15075_ (
);

OR2X2 _15360_ (
    .A(_4315_),
    .B(_4314_),
    .Y(_4316_)
);

FILL FILL_1__14815_ (
);

OR2X2 _16985_ (
    .A(_5900_),
    .B(_5915_),
    .Y(_5916_)
);

OR2X2 _16565_ (
    .A(_5502_),
    .B(_5501_),
    .Y(_5503_)
);

AND2X2 _16145_ (
    .A(_4214__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_5089_)
);

DFFSR _11280_ (
    .CLK(clk_bF$buf61),
    .D(_1389_[18]),
    .Q(\datapath_1.regfile_1.regOut[22] [18]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL_0__17641_ (
);

FILL FILL_0__17221_ (
);

FILL FILL395200x197600 (
);

FILL FILL108680x182780 (
);

OR2X2 _8487_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_23_)
);

FILL FILL492480x148200 (
);

OR2X2 _12485_ (
    .A(ALUOp[0]),
    .B(_2076_),
    .Y(ALUControl[2])
);

FILL FILL505400x148200 (
);

DFFSR _12065_ (
    .CLK(clk_bF$buf78),
    .D(_1785_[29]),
    .Q(\datapath_1.regfile_1.regOut[28] [29]),
    .R(rst_bF$buf110),
    .S(vdd)
);

FILL FILL414960x207480 (
);

FILL FILL_0__18846_ (
);

AND2X2 _18711_ (
    .A(_6323__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_7616_)
);

FILL FILL_0__18426_ (
);

FILL FILL_0__13981_ (
);

FILL FILL_0__13141_ (
);

FILL FILL131480x360620 (
);

FILL FILL_0__8527_ (
);

FILL FILL_1__9170_ (
);

FILL FILL285000x217360 (
);

FILL FILL427120x251940 (
);

FILL FILL_1__15773_ (
);

FILL FILL_0__14766_ (
);

OR2X2 _14631_ (
    .A(\datapath_1.rd1 [1]),
    .B(_3869__bF$buf1),
    .Y(_3807_)
);

AND2X2 _14211_ (
    .A(_3585_),
    .B(_3584_),
    .Y(\datapath_1.mux_wd3.dout [22])
);

FILL FILL253080x93860 (
);

FILL FILL249280x350740 (
);

FILL FILL285760x202540 (
);

FILL FILL_1__16978_ (
);

FILL FILL435480x365560 (
);

OR2X2 _15836_ (
    .A(_4783_),
    .B(_4784_),
    .Y(_4785_)
);

OR2X2 _15416_ (
    .A(_4356_),
    .B(_4371_),
    .Y(_4372_)
);

FILL FILL266760x360620 (
);

OR2X2 _10971_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_1299_)
);

FILL FILL_0__10266_ (
);

OR2X2 _10551_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_1079_)
);

DFFSR _10131_ (
    .CLK(clk_bF$buf7),
    .D(_795_[30]),
    .Q(\datapath_1.regfile_1.regOut[13] [30]),
    .R(rst_bF$buf48),
    .S(vdd)
);

FILL FILL5320x167960 (
);

FILL FILL_0__16912_ (
);

FILL FILL_0__19384_ (
);

FILL FILL201400x370500 (
);

FILL FILL_1__12478_ (
);

AND2X2 _11756_ (
    .A(_1702_),
    .B(_1701_),
    .Y(_1653_[24])
);

FILL FILL_0__9065_ (
);

AND2X2 _11336_ (
    .A(_1482_),
    .B(_1481_),
    .Y(_1455_[13])
);

FILL FILL_0__12832_ (
);

FILL FILL_0__12412_ (
);

FILL FILL277400x232180 (
);

FILL FILL290320x54340 (
);

FILL FILL60040x232180 (
);

OR2X2 _9904_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .B(_794__bF$buf1),
    .Y(_748_)
);

FILL FILL_1__8861_ (
);

FILL FILL319200x360620 (
);

FILL FILL163400x350740 (
);

FILL FILL329080x306280 (
);

AND2X2 _13902_ (
    .A(_3334_),
    .B(_3333_),
    .Y(\datapath_1.alu_1.ALUInA [28])
);

FILL FILL_0__13617_ (
);

FILL FILL505400x375440 (
);

FILL FILL209760x256880 (
);

FILL FILL_1__17096_ (
);

FILL FILL381520x153140 (
);

AND2X2 _16794_ (
    .A(_4158__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_5728_)
);

FILL FILL_0__16089_ (
);

OR2X2 _16374_ (
    .A(_5314_),
    .B(_5311_),
    .Y(_5315_)
);

FILL FILL_0__17870_ (
);

FILL FILL_0__17030_ (
);

BUFX2 BUFX2_insert580 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf59)
);

BUFX2 BUFX2_insert581 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf58)
);

BUFX2 BUFX2_insert582 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf57)
);

BUFX2 BUFX2_insert583 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf56)
);

FILL FILL456760x0 (
);

BUFX2 BUFX2_insert584 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf55)
);

AND2X2 _17999_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_6915_)
);

FILL FILL22800x59280 (
);

BUFX2 BUFX2_insert585 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf54)
);

INVX1 _17579_ (
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_6502_)
);

BUFX2 BUFX2_insert586 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf53)
);

OR2X2 _17159_ (
    .A(_6086_),
    .B(_6085_),
    .Y(_6087_)
);

BUFX2 BUFX2_insert587 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf52)
);

BUFX2 BUFX2_insert588 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf51)
);

BUFX2 BUFX2_insert589 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf50)
);

DFFSR _12294_ (
    .CLK(clk_bF$buf105),
    .D(_1917_[0]),
    .Q(\datapath_1.regfile_1.regOut[30] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

FILL FILL_1__19242_ (
);

FILL FILL499320x143260 (
);

AND2X2 _18940_ (
    .A(_6232__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_7842_)
);

FILL FILL_0__18235_ (
);

AND2X2 _18520_ (
    .A(_6232__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_7428_)
);

AND2X2 _18100_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_7015_)
);

FILL FILL85120x24700 (
);

FILL FILL_0__13790_ (
);

FILL FILL_0__13370_ (
);

FILL FILL399000x237120 (
);

FILL FILL_0__8756_ (
);

AND2X2 _10607_ (
    .A(_1116_),
    .B(_1115_),
    .Y(_1059_[28])
);

FILL FILL376960x138320 (
);

OR2X2 _13499_ (
    .A(ALUOut[3]),
    .B(_3079__bF$buf4),
    .Y(_3021_)
);

INVX1 _13079_ (
    .A(_2634_),
    .Y(\datapath_1.ALUResult [22])
);

AND2X2 _19305_ (
    .A(_6323__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_8201_)
);

DFFSR _14860_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[8]),
    .Q(_2_[8]),
    .R(rst_bF$buf61),
    .S(vdd)
);

FILL FILL_0__14575_ (
);

FILL FILL_0__14155_ (
);

AND2X2 _14440_ (
    .A(_3719_),
    .B(_3718_),
    .Y(_3672_[23])
);

AND2X2 _14020_ (
    .A(_3352__bF$buf0),
    .B(\datapath_1.PCJump [14]),
    .Y(_3437_)
);

AND2X2 _15645_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_4597_)
);

AND2X2 _15225_ (
    .A(_4141_),
    .B(_4171_),
    .Y(_4183_)
);

FILL FILL21280x69160 (
);

OR2X2 _10780_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(_1256__bF$buf2),
    .Y(_1192_)
);

DFFSR _10360_ (
    .CLK(clk_bF$buf21),
    .D(_927_[1]),
    .Q(\datapath_1.regfile_1.regOut[15] [1]),
    .R(rst_bF$buf90),
    .S(vdd)
);

FILL FILL142120x370500 (
);

FILL FILL172520x281580 (
);

FILL FILL133760x247000 (
);

FILL FILL256120x118560 (
);

FILL FILL50920x281580 (
);

FILL FILL_0__19193_ (
);

FILL FILL397480x296400 (
);

FILL FILL47880x232180 (
);

FILL FILL_0__9294_ (
);

OR2X2 _11985_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_1815_)
);

FILL FILL_1__18933_ (
);

OR2X2 _11565_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_1595_)
);

DFFSR _11145_ (
    .CLK(clk_bF$buf103),
    .D(_1323_[12]),
    .Q(\datapath_1.regfile_1.regOut[21] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

FILL FILL41800x256880 (
);

FILL FILL_0__17926_ (
);

FILL FILL_0__17506_ (
);

FILL FILL_0__12221_ (
);

FILL FILL345800x167960 (
);

AND2X2 _9713_ (
    .A(_660_),
    .B(_659_),
    .Y(_597_[31])
);

FILL FILL25080x69160 (
);

FILL FILL351120x335920 (
);

FILL FILL402040x29640 (
);

FILL FILL167960x266760 (
);

FILL FILL_0__13846_ (
);

FILL FILL_0__13426_ (
);

AND2X2 _13711_ (
    .A(_3084__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3189_)
);

FILL FILL_0__13006_ (
);

OR2X2 _16183_ (
    .A(_5119_),
    .B(_5126_),
    .Y(_5127_)
);

FILL FILL_1__9875_ (
);

FILL FILL_1__9455_ (
);

FILL FILL504640x143260 (
);

OR2X2 _14916_ (
    .A(\datapath_1.mux_pcsrc.dout [10]),
    .B(_4001__bF$buf3),
    .Y(_3957_)
);

OR2X2 _17388_ (
    .A(_6313_),
    .B(_6311_),
    .Y(_6314_)
);

FILL FILL_0__18884_ (
);

FILL FILL_0__18464_ (
);

FILL FILL_1__11558_ (
);

FILL FILL_0__8985_ (
);

OR2X2 _10836_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_1229_)
);

OR2X2 _10416_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_1009_)
);

DFFSR _19534_ (
    .CLK(clk_bF$buf45),
    .D(_8320_[11]),
    .Q(\datapath_1.regfile_1.regOut[0] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL_0__19249_ (
);

OR2X2 _19114_ (
    .A(_8009_),
    .B(_8012_),
    .Y(_8013_)
);

FILL FILL_0__14384_ (
);

FILL FILL138320x172900 (
);

FILL FILL20520x276640 (
);

FILL FILL343520x350740 (
);

FILL FILL151240x167960 (
);

FILL FILL326040x44460 (
);

FILL FILL258400x19760 (
);

FILL FILL_1__16596_ (
);

AND2X2 _15874_ (
    .A(_4200__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_4822_)
);

AND2X2 _15454_ (
    .A(_4183__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_4409_)
);

FILL FILL_0__15169_ (
);

OR2X2 _15034_ (
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_4023_)
);

FILL FILL146680x286520 (
);

FILL FILL_0__16530_ (
);

FILL FILL_0__16110_ (
);

OR2X2 _16659_ (
    .A(_5593_),
    .B(_5594_),
    .Y(_5595_)
);

OR2X2 _16239_ (
    .A(_5178_),
    .B(_5181_),
    .Y(_5182_)
);

DFFSR _11794_ (
    .CLK(clk_bF$buf53),
    .D(_1653_[16]),
    .Q(\datapath_1.regfile_1.regOut[26] [16]),
    .R(rst_bF$buf110),
    .S(vdd)
);

OR2X2 _11374_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .B(_1520__bF$buf3),
    .Y(_1508_)
);

FILL FILL_0__11089_ (
);

FILL FILL_0__17735_ (
);

OR2X2 _17600_ (
    .A(_6519_),
    .B(_6522_),
    .Y(_6523_)
);

FILL FILL_0__17315_ (
);

FILL FILL464360x29640 (
);

FILL FILL_0__12870_ (
);

FILL FILL_0__12030_ (
);

FILL FILL231800x217360 (
);

FILL FILL_1__10829_ (
);

FILL FILL132240x113620 (
);

FILL FILL216600x49400 (
);

OR2X2 _9942_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_773_)
);

OR2X2 _9522_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_553_)
);

INVX2 _9102_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .Y(_398_)
);

AOI21X1 _12999_ (
    .A(_2547_),
    .B(_2559_),
    .C(_2552_),
    .Y(_2560_)
);

OR2X2 _12579_ (
    .A(\control_1.next [2]),
    .B(_2145_),
    .Y(_2150_)
);

OR2X2 _12159_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_1911_)
);

FILL FILL_1__19107_ (
);

OR2X2 _18805_ (
    .A(_7694_),
    .B(_7708_),
    .Y(_7709_)
);

AND2X2 _13940_ (
    .A(_3347__bF$buf2),
    .B(\aluControl_1.inst [3]),
    .Y(_3368_)
);

FILL FILL_0__13655_ (
);

OR2X2 _13520_ (
    .A(ALUOut[10]),
    .B(_3079__bF$buf0),
    .Y(_3035_)
);

FILL FILL_0_BUFX2_insert225 (
);

XOR2X1 _13100_ (
    .A(_2274_),
    .B(_2601_),
    .Y(_2654_)
);

FILL FILL_0_BUFX2_insert227 (
);

FILL FILL_0_BUFX2_insert229 (
);

BUFX2 BUFX2_insert1140 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf4 )
);

BUFX2 BUFX2_insert1141 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf3 )
);

BUFX2 BUFX2_insert1142 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf2 )
);

BUFX2 BUFX2_insert1143 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf1 )
);

BUFX2 BUFX2_insert1144 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf0 )
);

BUFX2 BUFX2_insert1145 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf4 )
);

FILL FILL322240x370500 (
);

BUFX2 BUFX2_insert1146 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf3 )
);

BUFX2 BUFX2_insert1147 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf2 )
);

BUFX2 BUFX2_insert1148 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf1 )
);

FILL FILL_1__15447_ (
);

FILL FILL113240x64220 (
);

BUFX2 BUFX2_insert1149 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf0 )
);

FILL FILL_1__10582_ (
);

DFFSR _14725_ (
    .CLK(clk_bF$buf58),
    .D(_3804_[2]),
    .Q(\datapath_1.a [2]),
    .R(rst_bF$buf15),
    .S(vdd)
);

AND2X2 _14305_ (
    .A(_3649_),
    .B(_3648_),
    .Y(_3606_[21])
);

BUFX2 BUFX2_insert960 (
    .A(_6211_),
    .Y(_6211__bF$buf0)
);

BUFX2 BUFX2_insert961 (
    .A(_1916_),
    .Y(_1916__bF$buf4)
);

BUFX2 BUFX2_insert962 (
    .A(_1916_),
    .Y(_1916__bF$buf3)
);

BUFX2 BUFX2_insert963 (
    .A(_1916_),
    .Y(_1916__bF$buf2)
);

BUFX2 BUFX2_insert964 (
    .A(_1916_),
    .Y(_1916__bF$buf1)
);

BUFX2 BUFX2_insert965 (
    .A(_1916_),
    .Y(_1916__bF$buf0)
);

BUFX2 BUFX2_insert966 (
    .A(_4197_),
    .Y(_4197__bF$buf4)
);

AND2X2 _17197_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_6125_)
);

BUFX2 BUFX2_insert967 (
    .A(_4197_),
    .Y(_4197__bF$buf3)
);

FILL FILL392920x158080 (
);

BUFX2 BUFX2_insert968 (
    .A(_4197_),
    .Y(_4197__bF$buf2)
);

BUFX2 BUFX2_insert969 (
    .A(_4197_),
    .Y(_4197__bF$buf1)
);

FILL FILL_1__19280_ (
);

FILL FILL197600x118560 (
);

FILL FILL_0__18693_ (
);

FILL FILL388360x44460 (
);

FILL FILL_0__8794_ (
);

DFFSR _10645_ (
    .CLK(clk_bF$buf110),
    .D(_1059_[28]),
    .Q(\datapath_1.regfile_1.regOut[17] [28]),
    .R(rst_bF$buf74),
    .S(vdd)
);

OR2X2 _10225_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .B(_926__bF$buf3),
    .Y(_922_)
);

FILL FILL478800x83980 (
);

FILL FILL_0__11721_ (
);

FILL FILL_0__19478_ (
);

FILL FILL_0__19058_ (
);

AND2X2 _19343_ (
    .A(_6297__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_8239_)
);

FILL FILL_0__14193_ (
);

FILL FILL298680x311220 (
);

FILL FILL_0__9579_ (
);

FILL FILL288040x271700 (
);

FILL FILL_1__13513_ (
);

FILL FILL_0__15398_ (
);

AND2X2 _15683_ (
    .A(_4160__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_4634_)
);

OR2X2 _15263_ (
    .A(_4206_),
    .B(_4220_),
    .Y(_4221_)
);

FILL FILL428640x133380 (
);

FILL FILL411160x217360 (
);

OR2X2 _16888_ (
    .A(_5805_),
    .B(_5820_),
    .Y(_5821_)
);

AND2X2 _16468_ (
    .A(_4175__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_5407_)
);

AND2X2 _16048_ (
    .A(_4151__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_4994_)
);

AND2X2 _11183_ (
    .A(_1400_),
    .B(_1399_),
    .Y(_1389_[5])
);

FILL FILL28120x237120 (
);

FILL FILL_0__17964_ (
);

FILL FILL_0__17544_ (
);

FILL FILL500840x266760 (
);

OR2X2 _9751_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .B(_728__bF$buf3),
    .Y(_666_)
);

DFFSR _9331_ (
    .CLK(clk_bF$buf51),
    .D(_399_[4]),
    .Q(\datapath_1.regfile_1.regOut[7] [4]),
    .R(rst_bF$buf83),
    .S(vdd)
);

OR2X2 _12388_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_2048__bF$buf1),
    .Y(_2024_)
);

OR2X2 _18614_ (
    .A(_7519_),
    .B(_7520_),
    .Y(_7521_)
);

FILL FILL_0__18329_ (
);

FILL FILL_0__13464_ (
);

FILL FILL_0__13044_ (
);

FILL FILL_0__14669_ (
);

OR2X2 _14954_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [23]),
    .Y(_3982_)
);

OR2X2 _14534_ (
    .A(IRWrite_bF$buf0),
    .B(\datapath_1.PCJump [14]),
    .Y(_3762_)
);

AND2X2 _14114_ (
    .A(_3344__bF$buf1),
    .B(gnd),
    .Y(_3517_)
);

FILL FILL_0__15610_ (
);

FILL FILL_0__18082_ (
);

FILL FILL407360x153140 (
);

FILL FILL196080x14820 (
);

AND2X2 _15739_ (
    .A(_4195__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_4689_)
);

OR2X2 _15319_ (
    .A(_4272_),
    .B(_4275_),
    .Y(_4276_)
);

FILL FILL206720x360620 (
);

AND2X2 _10874_ (
    .A(_1254_),
    .B(_1253_),
    .Y(_1191_[31])
);

AND2X2 _10454_ (
    .A(_1034_),
    .B(_1033_),
    .Y(_993_[20])
);

FILL FILL_0__10169_ (
);

FILL FILL_1__17402_ (
);

AND2X2 _10034_ (
    .A(_814_),
    .B(_813_),
    .Y(_795_[9])
);

FILL FILL_0__11950_ (
);

FILL FILL_0__11110_ (
);

FILL FILL_0__19287_ (
);

OR2X2 _19152_ (
    .A(_8050_),
    .B(_8049_),
    .Y(_8051_)
);

OR2X2 _8602_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .B(_134__bF$buf2),
    .Y(_80_)
);

FILL FILL_0__9388_ (
);

FILL FILL_1__18607_ (
);

DFFSR _11659_ (
    .CLK(clk_bF$buf0),
    .D(_1587_[10]),
    .Q(\datapath_1.regfile_1.regOut[25] [10]),
    .R(rst_bF$buf37),
    .S(vdd)
);

OR2X2 _11239_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_1454__bF$buf4),
    .Y(_1438_)
);

FILL FILL_0__12735_ (
);

NAND2X1 _12600_ (
    .A(_2164_),
    .B(_2161_),
    .Y(_2165_)
);

FILL FILL57000x88920 (
);

OR2X2 _15492_ (
    .A(_4444_),
    .B(_4445_),
    .Y(_4446_)
);

NOR2X1 _15072_ (
    .A(_4054_),
    .B(\datapath_1.a3 [0]),
    .Y(_4059_)
);

OR2X2 _9807_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_703_)
);

FILL FILL37240x355680 (
);

FILL FILL_1__14947_ (
);

AND2X2 _13805_ (
    .A(_3089__bF$buf1),
    .B(gnd),
    .Y(_3270_)
);

OR2X2 _16697_ (
    .A(_5601_),
    .B(_5632_),
    .Y(_5633_)
);

AND2X2 _16277_ (
    .A(_4210__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_5219_)
);

FILL FILL_1__18360_ (
);

FILL FILL_0__17353_ (
);

FILL FILL130720x306280 (
);

DFFSR _9980_ (
    .CLK(clk_bF$buf52),
    .D(_729_[8]),
    .Q(\datapath_1.regfile_1.regOut[12] [8]),
    .R(rst_bF$buf0),
    .S(vdd)
);

AND2X2 _9560_ (
    .A(_578_),
    .B(_577_),
    .Y(_531_[23])
);

AND2X2 _9140_ (
    .A(_358_),
    .B(_357_),
    .Y(_333_[12])
);

OR2X2 _12197_ (
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .Y(_1981_)
);

FILL FILL_0__10801_ (
);

FILL FILL_0__18978_ (
);

FILL FILL_0_BUFX2_insert600 (
);

FILL FILL_0__18558_ (
);

OR2X2 _18843_ (
    .A(_7745_),
    .B(_7744_),
    .Y(_7746_)
);

FILL FILL_0_BUFX2_insert601 (
);

AND2X2 _18423_ (
    .A(_6255__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_7333_)
);

AND2X2 _18003_ (
    .A(_6315__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_6919_)
);

FILL FILL_0_BUFX2_insert603 (
);

FILL FILL_0__13693_ (
);

FILL FILL_0__13273_ (
);

FILL FILL_0_BUFX2_insert605 (
);

FILL FILL_0_BUFX2_insert607 (
);

FILL FILL_0_BUFX2_insert609 (
);

FILL FILL504640x306280 (
);

FILL FILL_1__15065_ (
);

OR2X2 _19208_ (
    .A(_8104_),
    .B(_8105_),
    .Y(_8106_)
);

FILL FILL_0__14898_ (
);

FILL FILL414960x54340 (
);

OR2X2 _14763_ (
    .A(\datapath_1.rd2 [2]),
    .B(_3935__bF$buf2),
    .Y(_3875_)
);

FILL FILL_0__14058_ (
);

DFFSR _14343_ (
    .CLK(clk_bF$buf12),
    .D(_3606_[7]),
    .Q(ALUOut[7]),
    .R(rst_bF$buf91),
    .S(vdd)
);

FILL FILL278160x158080 (
);

FILL FILL10640x79040 (
);

OR2X2 _15968_ (
    .A(_4911_),
    .B(_4914_),
    .Y(_4915_)
);

FILL FILL411160x69160 (
);

AND2X2 _15548_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_4501_)
);

NAND3X1 _15128_ (
    .A(_4031_),
    .B(_4054_),
    .C(_4017_),
    .Y(_4104_)
);

OR2X2 _10683_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_1147_)
);

FILL FILL270560x123500 (
);

INVX2 _10263_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .Y(_992_)
);

FILL FILL_0__16204_ (
);

OR2X2 _19381_ (
    .A(_8271_),
    .B(_8275_),
    .Y(_8276_)
);

DFFSR _8831_ (
    .CLK(clk_bF$buf100),
    .D(_135_[20]),
    .Q(\datapath_1.regfile_1.regOut[3] [20]),
    .R(rst_bF$buf68),
    .S(vdd)
);

BUFX2 _8411_ (
    .A(_1_[19]),
    .Y(memoryAddress[19])
);

AND2X2 _11888_ (
    .A(_1770_),
    .B(_1769_),
    .Y(_1719_[25])
);

FILL FILL_0__9197_ (
);

AND2X2 _11468_ (
    .A(_1550_),
    .B(_1549_),
    .Y(_1521_[14])
);

AND2X2 _11048_ (
    .A(_1330_),
    .B(_1329_),
    .Y(_1323_[3])
);

FILL FILL_0__17829_ (
);

FILL FILL_0__17409_ (
);

FILL FILL126920x83980 (
);

FILL FILL78280x59280 (
);

FILL FILL_0__12964_ (
);

FILL FILL_0__12544_ (
);

FILL FILL240160x59280 (
);

DFFSR _9616_ (
    .CLK(clk_bF$buf27),
    .D(_531_[31]),
    .Q(\datapath_1.regfile_1.regOut[9] [31]),
    .R(rst_bF$buf28),
    .S(vdd)
);

FILL FILL_1__8993_ (
);

FILL FILL88160x123500 (
);

FILL FILL_1__14756_ (
);

FILL FILL30400x281580 (
);

OR2X2 _13614_ (
    .A(_3104_),
    .B(_3105_),
    .Y(_3106_)
);

OR2X2 _16086_ (
    .A(_5030_),
    .B(_5029_),
    .Y(_5031_)
);

FILL FILL38760x14820 (
);

FILL FILL_0__17582_ (
);

FILL FILL267520x59280 (
);

FILL FILL70680x4940 (
);

OR2X2 _14819_ (
    .A(vdd),
    .B(_2_[21]),
    .Y(_3912_)
);

FILL FILL_1__16902_ (
);

FILL FILL459040x19760 (
);

FILL FILL_1__19374_ (
);

FILL FILL_0__10610_ (
);

OR2X2 _18652_ (
    .A(_7557_),
    .B(_7554_),
    .Y(_7558_)
);

FILL FILL_0__18367_ (
);

FILL FILL354160x321100 (
);

AND2X2 _18232_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_7145_)
);

FILL FILL15960x88920 (
);

FILL FILL_0__8888_ (
);

AND2X2 _10739_ (
    .A(_1184_),
    .B(_1183_),
    .Y(_1125_[29])
);

AND2X2 _10319_ (
    .A(_964_),
    .B(_963_),
    .Y(_927_[18])
);

FILL FILL_1__12402_ (
);

OR2X2 _19437_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8327_)
);

FILL FILL93480x133380 (
);

NOR2X1 _19017_ (
    .A(_6310__bF$buf3),
    .B(_7917_),
    .Y(_7918_)
);

DFFSR _14992_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[11]),
    .Q(\datapath_1.mux_iord.din0 [11]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL_0__14287_ (
);

AND2X2 _14572_ (
    .A(_3787_),
    .B(_3786_),
    .Y(_3738_[24])
);

OR2X2 _14152_ (
    .A(MemToReg_bF$buf3),
    .B(ALUOut[3]),
    .Y(_3546_)
);

FILL FILL466640x237120 (
);

FILL FILL22040x83980 (
);

FILL FILL388360x340860 (
);

AND2X2 _15777_ (
    .A(_4203__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_4727_)
);

OR2X2 _15357_ (
    .A(_4312_),
    .B(_4311_),
    .Y(_4313_)
);

FILL FILL_1__17860_ (
);

DFFSR _10492_ (
    .CLK(clk_bF$buf82),
    .D(_993_[4]),
    .Q(\datapath_1.regfile_1.regOut[16] [4]),
    .R(rst_bF$buf94),
    .S(vdd)
);

OR2X2 _10072_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .B(_860__bF$buf0),
    .Y(_840_)
);

FILL FILL_0__16853_ (
);

FILL FILL_0__16433_ (
);

FILL FILL_0__16013_ (
);

AND2X2 _19190_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_8088_)
);

OR2X2 _8640_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_105_)
);

FILL FILL109440x370500 (
);

FILL FILL319200x54340 (
);

OR2X2 _11697_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_1663_)
);

FILL FILL_1__18225_ (
);

DFFSR _11277_ (
    .CLK(clk_bF$buf54),
    .D(_1389_[15]),
    .Q(\datapath_1.regfile_1.regOut[22] [15]),
    .R(rst_bF$buf24),
    .S(vdd)
);

AND2X2 _17923_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_6841_)
);

OR2X2 _17503_ (
    .A(_6426_),
    .B(_6423_),
    .Y(_6427_)
);

FILL FILL_0__12773_ (
);

FILL FILL505400x261820 (
);

FILL FILL_0__12353_ (
);

FILL FILL430160x39520 (
);

DFFSR _9845_ (
    .CLK(clk_bF$buf18),
    .D(_663_[2]),
    .Q(\datapath_1.regfile_1.regOut[11] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _9425_ (
    .A(_508_),
    .B(_507_),
    .Y(_465_[21])
);

FILL FILL23560x128440 (
);

AND2X2 _9005_ (
    .A(_288_),
    .B(_287_),
    .Y(_267_[10])
);

FILL FILL262960x14820 (
);

FILL FILL285000x330980 (
);

OR2X2 _18708_ (
    .A(_7582_),
    .B(_7613_),
    .Y(_7614_)
);

FILL FILL276640x207480 (
);

OR2X2 _13843_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [9]),
    .Y(_3295_)
);

FILL FILL_0__13558_ (
);

FILL FILL_0__13138_ (
);

OR2X2 _13423_ (
    .A(_2957_),
    .B(_2387__bF$buf0),
    .Y(_2958_)
);

FILL FILL350360x54340 (
);

OR2X2 _13003_ (
    .A(_2157__bF$buf2),
    .B(_2562_),
    .Y(_2563_)
);

FILL FILL177080x103740 (
);

FILL FILL353400x172900 (
);

FILL FILL450680x123500 (
);

OR2X2 _14628_ (
    .A(\datapath_1.rd1 [0]),
    .B(_3869__bF$buf0),
    .Y(_3805_)
);

AND2X2 _14208_ (
    .A(_3583_),
    .B(_3582_),
    .Y(\datapath_1.mux_wd3.dout [21])
);

FILL FILL335920x345800 (
);

FILL FILL_0__15704_ (
);

FILL FILL338200x232180 (
);

FILL FILL52440x9880 (
);

AND2X2 _18881_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_7784_)
);

FILL FILL_0__18176_ (
);

AND2X2 _18461_ (
    .A(_6315__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_7370_)
);

INVX1 _18041_ (
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_6957_)
);

FILL FILL330600x24700 (
);

OR2X2 _10968_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_1297_)
);

OR2X2 _10548_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_1077_)
);

DFFSR _10128_ (
    .CLK(clk_bF$buf36),
    .D(_795_[27]),
    .Q(\datapath_1.regfile_1.regOut[13] [27]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL_1__12631_ (
);

FILL FILL_0__16909_ (
);

FILL FILL_0__11624_ (
);

AND2X2 _19246_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_8143_)
);

FILL FILL247000x113620 (
);

FILL FILL_0__14096_ (
);

OR2X2 _14381_ (
    .A(vdd),
    .B(\datapath_1.Data [4]),
    .Y(_3680_)
);

FILL FILL407360x316160 (
);

FILL FILL421040x93860 (
);

FILL FILL390640x44460 (
);

FILL FILL219640x148200 (
);

FILL FILL_0__12829_ (
);

AND2X2 _15586_ (
    .A(_4160__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_4539_)
);

NOR3X1 _15166_ (
    .A(_4125_),
    .B(_4054_),
    .C(_4010_),
    .Y(\datapath_1.regfile_1.regEn [30])
);

FILL FILL336680x291460 (
);

FILL FILL255360x227240 (
);

FILL FILL_0__16662_ (
);

FILL FILL492480x39520 (
);

FILL FILL88160x83980 (
);

FILL FILL395200x108680 (
);

FILL FILL482600x113620 (
);

FILL FILL_1__18874_ (
);

OR2X2 _11086_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .B(_1388__bF$buf1),
    .Y(_1356_)
);

FILL FILL_0__17447_ (
);

OR2X2 _17732_ (
    .A(_6637_),
    .B(_6652_),
    .Y(_6653_)
);

FILL FILL_0__17027_ (
);

AND2X2 _17312_ (
    .A(_6205_),
    .B(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_6238_)
);

FILL FILL_0__12582_ (
);

FILL FILL_0__12162_ (
);

FILL FILL86640x316160 (
);

FILL FILL36480x167960 (
);

OR2X2 _9654_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_621_)
);

OR2X2 _9234_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_401_)
);

FILL FILL76000x276640 (
);

FILL FILL_1__11902_ (
);

FILL FILL72960x340860 (
);

AND2X2 _18937_ (
    .A(_6272__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_7839_)
);

AND2X2 _18517_ (
    .A(_6216__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_7425_)
);

FILL FILL259160x335920 (
);

FILL FILL_0__13787_ (
);

OR2X2 _13652_ (
    .A(_3138_),
    .B(_3137_),
    .Y(_3139_)
);

INVX1 _13232_ (
    .A(_2778_),
    .Y(\datapath_1.ALUResult [13])
);

FILL FILL494760x148200 (
);

FILL FILL_1__15579_ (
);

FILL FILL230280x326040 (
);

DFFSR _14857_ (
    .CLK(clk_bF$buf15),
    .D(_3870_[5]),
    .Q(_2_[5]),
    .R(rst_bF$buf53),
    .S(vdd)
);

AND2X2 _14437_ (
    .A(_3717_),
    .B(_3716_),
    .Y(_3672_[22])
);

AND2X2 _14017_ (
    .A(_3347__bF$buf1),
    .B(\datapath_1.PCJump [16]),
    .Y(_3434_)
);

FILL FILL_0_CLKBUF1_insert211 (
);

FILL FILL_0__15933_ (
);

FILL FILL_0_CLKBUF1_insert213 (
);

FILL FILL_0__15513_ (
);

FILL FILL_0_CLKBUF1_insert215 (
);

FILL FILL_0_CLKBUF1_insert217 (
);

FILL FILL_0_CLKBUF1_insert218 (
);

FILL FILL_0_CLKBUF1_insert219 (
);

OR2X2 _18690_ (
    .A(_7592_),
    .B(_7595_),
    .Y(_7596_)
);

OR2X2 _18270_ (
    .A(_7181_),
    .B(_7174_),
    .Y(_7182_)
);

FILL FILL133760x360620 (
);

FILL FILL114760x197600 (
);

FILL FILL429400x251940 (
);

FILL FILL57000x222300 (
);

DFFSR _10777_ (
    .CLK(clk_bF$buf100),
    .D(_1125_[31]),
    .Q(\datapath_1.regfile_1.regOut[18] [31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL_1__17725_ (
);

OR2X2 _10357_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .B(_992__bF$buf0),
    .Y(_990_)
);

FILL FILL_1__12020_ (
);

FILL FILL_0__16718_ (
);

FILL FILL_0__11853_ (
);

FILL FILL_0__11433_ (
);

OR2X2 _19475_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_8352_)
);

OR2X2 _19055_ (
    .A(_7953_),
    .B(_7954_),
    .Y(_7955_)
);

AND2X2 _14190_ (
    .A(_3571_),
    .B(_3570_),
    .Y(\datapath_1.mux_wd3.dout [15])
);

OR2X2 _8925_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_255_)
);

OR2X2 _8505_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_35_)
);

FILL FILL211280x34580 (
);

FILL FILL_1_BUFX2_insert531 (
);

NOR2X1 _12923_ (
    .A(_2487_),
    .B(_2353_),
    .Y(_2488_)
);

FILL FILL_0__12638_ (
);

INVX1 _12503_ (
    .A(\control_1.reg_state.dout [3]),
    .Y(_2100_)
);

FILL FILL_1_BUFX2_insert533 (
);

FILL FILL51680x360620 (
);

FILL FILL7600x167960 (
);

OR2X2 _15395_ (
    .A(_4349_),
    .B(_4350_),
    .Y(_4351_)
);

FILL FILL318440x19760 (
);

FILL FILL_0__16051_ (
);

FILL FILL400520x108680 (
);

OR2X2 _13708_ (
    .A(_3186_),
    .B(_3185_),
    .Y(_3187_)
);

FILL FILL285760x276640 (
);

FILL FILL373920x98800 (
);

AND2X2 _17961_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_6878_)
);

FILL FILL_0__17676_ (
);

AND2X2 _17541_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_6464_)
);

AND2X2 _17121_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_6050_)
);

FILL FILL_0__12391_ (
);

OR2X2 _9883_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_794__bF$buf4),
    .Y(_734_)
);

DFFSR _9463_ (
    .CLK(clk_bF$buf18),
    .D(_465_[7]),
    .Q(\datapath_1.regfile_1.regOut[8] [7]),
    .R(rst_bF$buf3),
    .S(vdd)
);

OR2X2 _9043_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .B(_332__bF$buf4),
    .Y(_314_)
);

FILL FILL_1__11711_ (
);

FILL FILL101840x39520 (
);

FILL FILL_1__19048_ (
);

FILL FILL_0__10704_ (
);

AND2X2 _18746_ (
    .A(_6232__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [21]),
    .Y(_7651_)
);

NOR2X1 _18326_ (
    .A(_6310__bF$buf0),
    .B(_7236_),
    .Y(_7237_)
);

AND2X2 _13881_ (
    .A(_3320_),
    .B(_3319_),
    .Y(\datapath_1.alu_1.ALUInA [21])
);

FILL FILL_0__13176_ (
);

AND2X2 _13461_ (
    .A(_2993_),
    .B(_2889_),
    .Y(_2994_)
);

AND2X2 _13041_ (
    .A(_2598_),
    .B(_2589_),
    .Y(_2599_)
);

FILL FILL88160x0 (
);

FILL FILL_0__9503_ (
);

OR2X2 _14666_ (
    .A(vdd),
    .B(\datapath_1.a [13]),
    .Y(_3830_)
);

OR2X2 _14246_ (
    .A(vdd),
    .B(ALUOut[2]),
    .Y(_3610_)
);

FILL FILL57760x217360 (
);

FILL FILL169480x19760 (
);

FILL FILL364800x177840 (
);

FILL FILL_0__15322_ (
);

BUFX2 BUFX2_insert0 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf4 )
);

BUFX2 BUFX2_insert1 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf3 )
);

BUFX2 BUFX2_insert2 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf2 )
);

BUFX2 BUFX2_insert3 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf1 )
);

BUFX2 BUFX2_insert4 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf0 )
);

BUFX2 BUFX2_insert5 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf4 )
);

BUFX2 BUFX2_insert6 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf3 )
);

FILL FILL105640x39520 (
);

BUFX2 BUFX2_insert7 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf2 )
);

BUFX2 BUFX2_insert8 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf1 )
);

BUFX2 BUFX2_insert9 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf0 )
);

FILL FILL64600x187720 (
);

FILL FILL204440x182780 (
);

FILL FILL_1__17954_ (
);

AND2X2 _10586_ (
    .A(_1102_),
    .B(_1101_),
    .Y(_1059_[21])
);

AND2X2 _10166_ (
    .A(_882_),
    .B(_881_),
    .Y(_861_[10])
);

FILL FILL397480x207480 (
);

FILL FILL_0__16947_ (
);

FILL FILL_0__16527_ (
);

AND2X2 _16812_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_5746_)
);

FILL FILL264480x296400 (
);

FILL FILL_0__11242_ (
);

AND2X2 _19284_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_8181_)
);

FILL FILL85120x98800 (
);

OR2X2 _8734_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .B(_200__bF$buf3),
    .Y(_148_)
);

FILL FILL_1__18739_ (
);

FILL FILL_1__13454_ (
);

FILL FILL_1__13034_ (
);

NAND2X1 _12732_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(_2296_),
    .Y(_2297_)
);

DFFSR _12312_ (
    .CLK(clk_bF$buf52),
    .D(_1917_[18]),
    .Q(\datapath_1.regfile_1.regOut[30] [18]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL_0__12027_ (
);

FILL FILL144400x370500 (
);

FILL FILL484880x34580 (
);

OR2X2 _9939_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_771_)
);

OR2X2 _9519_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_551_)
);

FILL FILL_1__8896_ (
);

FILL FILL_0__16280_ (
);

FILL FILL39520x192660 (
);

OR2X2 _13937_ (
    .A(_3365_),
    .B(_3364_),
    .Y(_3366_)
);

OR2X2 _13517_ (
    .A(ALUOut[9]),
    .B(_3079__bF$buf3),
    .Y(_3033_)
);

FILL FILL161120x286520 (
);

FILL FILL_0__17485_ (
);

AND2X2 _17770_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_6690_)
);

FILL FILL_0__17065_ (
);

NOR2X1 _17350_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(\datapath_1.PCJump [26]),
    .Y(_6276_)
);

FILL FILL250040x19760 (
);

FILL FILL338960x49400 (
);

AND2X2 _9692_ (
    .A(_646_),
    .B(_645_),
    .Y(_597_[24])
);

AND2X2 _9272_ (
    .A(_426_),
    .B(_425_),
    .Y(_399_[13])
);

FILL FILL_1__11100_ (
);

FILL FILL_0__10933_ (
);

AND2X2 _18975_ (
    .A(_6221__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_7876_)
);

AND2X2 _18555_ (
    .A(_6326__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_7463_)
);

OR2X2 _18135_ (
    .A(_7048_),
    .B(_7047_),
    .Y(_7049_)
);

AND2X2 _13690_ (
    .A(_3084__bF$buf1),
    .B(\datapath_1.PCJump [14]),
    .Y(_3171_)
);

OAI21X1 _13270_ (
    .A(_2500_),
    .B(_2800_),
    .C(_2813_),
    .Y(_2814_)
);

FILL FILL_0__19211_ (
);

FILL FILL_0__11718_ (
);

FILL FILL_0__9312_ (
);

OR2X2 _14895_ (
    .A(\datapath_1.mux_pcsrc.dout [3]),
    .B(_4001__bF$buf1),
    .Y(_3943_)
);

DFFSR _14475_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[10]),
    .Q(\datapath_1.Data [10]),
    .R(rst_bF$buf85),
    .S(vdd)
);

AND2X2 _14055_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3467_)
);

FILL FILL161880x9880 (
);

FILL FILL_0__15971_ (
);

FILL FILL_0__15551_ (
);

FILL FILL_0__15131_ (
);

FILL FILL15960x306280 (
);

FILL FILL328320x340860 (
);

FILL FILL273600x311220 (
);

OR2X2 _10395_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_995_)
);

FILL FILL_1__17343_ (
);

FILL FILL409640x88920 (
);

FILL FILL309320x177840 (
);

AND2X2 _16621_ (
    .A(_4175__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_5558_)
);

OR2X2 _16201_ (
    .A(_5143_),
    .B(_5136_),
    .Y(_5144_)
);

FILL FILL_0__11471_ (
);

FILL FILL22800x276640 (
);

FILL FILL_0__11051_ (
);

FILL FILL345800x350740 (
);

FILL FILL110200x54340 (
);

FILL FILL160360x9880 (
);

AND2X2 _19093_ (
    .A(_6297__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_7993_)
);

FILL FILL237880x123500 (
);

DFFSR _8963_ (
    .CLK(clk_bF$buf74),
    .D(_201_[23]),
    .Q(\datapath_1.regfile_1.regOut[4] [23]),
    .R(rst_bF$buf47),
    .S(vdd)
);

AND2X2 _8543_ (
    .A(_60_),
    .B(_59_),
    .Y(_3_[28])
);

FILL FILL_1__13683_ (
);

AND2X2 _17826_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_6745_)
);

OR2X2 _17406_ (
    .A(_6320_),
    .B(_6331_),
    .Y(_6332_)
);

FILL FILL_1_BUFX2_insert911 (
);

FILL FILL_0__12676_ (
);

INVX1 _12961_ (
    .A(_2157__bF$buf0),
    .Y(_2524_)
);

AND2X2 _12541_ (
    .A(_2108_),
    .B(_2110_),
    .Y(_2130_)
);

FILL FILL_1_BUFX2_insert913 (
);

FILL FILL111720x163020 (
);

OR2X2 _12121_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .B(_1916__bF$buf1),
    .Y(_1886_)
);

OR2X2 _9748_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_728__bF$buf0),
    .Y(_664_)
);

DFFSR _9328_ (
    .CLK(clk_bF$buf93),
    .D(_399_[1]),
    .Q(\datapath_1.regfile_1.regOut[7] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL_1__14888_ (
);

FILL FILL199880x103740 (
);

FILL FILL216600x207480 (
);

FILL FILL58520x172900 (
);

AND2X2 _13746_ (
    .A(_3084__bF$buf2),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_3219_)
);

FILL FILL184680x365560 (
);

AOI22X1 _13326_ (
    .A(_2202_),
    .B(_2504_),
    .C(_2548_),
    .D(_2866_),
    .Y(_2867_)
);

FILL FILL_0__14822_ (
);

FILL FILL_0__17294_ (
);

FILL FILL134520x113620 (
);

DFFSR _9081_ (
    .CLK(clk_bF$buf113),
    .D(_267_[12]),
    .Q(\datapath_1.regfile_1.regOut[5] [12]),
    .R(rst_bF$buf102),
    .S(vdd)
);

FILL FILL_0__10742_ (
);

FILL FILL_0__10322_ (
);

FILL FILL307040x360620 (
);

AND2X2 _18784_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_7688_)
);

FILL FILL_0__18499_ (
);

OR2X2 _18364_ (
    .A(_7274_),
    .B(_7273_),
    .Y(_7275_)
);

FILL FILL343520x64220 (
);

FILL FILL_0__19440_ (
);

FILL FILL_1__17819_ (
);

FILL FILL352640x103740 (
);

FILL FILL_0__9541_ (
);

OR2X2 _11812_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(_1784__bF$buf2),
    .Y(_1720_)
);

FILL FILL_0__9121_ (
);

FILL FILL_0__11107_ (
);

FILL FILL165680x311220 (
);

OR2X2 _19149_ (
    .A(_8047_),
    .B(_8045_),
    .Y(_8048_)
);

AND2X2 _14284_ (
    .A(_3635_),
    .B(_3634_),
    .Y(_3606_[14])
);

FILL FILL_0__15780_ (
);

FILL FILL_1__13319_ (
);

OR2X2 _15489_ (
    .A(_4439_),
    .B(_4442_),
    .Y(_4443_)
);

AND2X2 _15069_ (
    .A(_4056_),
    .B(_4047_),
    .Y(_4057_)
);

FILL FILL_1__17992_ (
);

FILL FILL472720x365560 (
);

FILL FILL_0__16565_ (
);

AND2X2 _16850_ (
    .A(_4223__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_5783_)
);

FILL FILL_0__16145_ (
);

OR2X2 _16430_ (
    .A(_5369_),
    .B(_5368_),
    .Y(_5370_)
);

AND2X2 _16010_ (
    .A(_4214__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_4956_)
);

FILL FILL50160x187720 (
);

FILL FILL_1__9702_ (
);

FILL FILL478040x83980 (
);

FILL FILL459040x276640 (
);

FILL FILL274360x49400 (
);

OR2X2 _8772_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_173_)
);

FILL FILL199880x330980 (
);

FILL FILL_1__13072_ (
);

OR2X2 _17635_ (
    .A(_6543_),
    .B(_6556_),
    .Y(_6557_)
);

AND2X2 _17215_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_6142_)
);

NAND2X1 _12770_ (
    .A(_2331_),
    .B(_2334_),
    .Y(_2335_)
);

FILL FILL_0__12485_ (
);

AND2X2 _12350_ (
    .A(_1998_),
    .B(_1997_),
    .Y(_1983_[7])
);

FILL FILL_0__18711_ (
);

FILL FILL413440x217360 (
);

DFFSR _9977_ (
    .CLK(clk_bF$buf36),
    .D(_729_[5]),
    .Q(\datapath_1.regfile_1.regOut[12] [5]),
    .R(rst_bF$buf78),
    .S(vdd)
);

AND2X2 _9557_ (
    .A(_576_),
    .B(_575_),
    .Y(_531_[22])
);

AND2X2 _9137_ (
    .A(_356_),
    .B(_355_),
    .Y(_333_[11])
);

FILL FILL_1__14697_ (
);

FILL FILL_0_BUFX2_insert570 (
);

FILL FILL436240x301340 (
);

FILL FILL_0_BUFX2_insert572 (
);

FILL FILL_0_BUFX2_insert573 (
);

AND2X2 _13975_ (
    .A(_3347__bF$buf1),
    .B(\datapath_1.PCJump [10]),
    .Y(_3398_)
);

FILL FILL_0_BUFX2_insert574 (
);

OR2X2 _13555_ (
    .A(IorD_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [22]),
    .Y(_3058_)
);

FILL FILL_0_BUFX2_insert575 (
);

OR2X2 _13135_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2687_)
);

FILL FILL_0_BUFX2_insert576 (
);

FILL FILL_0_BUFX2_insert578 (
);

FILL FILL164920x9880 (
);

FILL FILL_0__14631_ (
);

FILL FILL16720x261820 (
);

FILL FILL_1__16843_ (
);

FILL FILL_1__16423_ (
);

FILL FILL_0__15416_ (
);

AND2X2 _15701_ (
    .A(_4189__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_4652_)
);

FILL FILL327560x59280 (
);

FILL FILL_0__10551_ (
);

OR2X2 _18593_ (
    .A(_7499_),
    .B(_7498_),
    .Y(_7500_)
);

OR2X2 _18173_ (
    .A(_7086_),
    .B(_7085_),
    .Y(_7087_)
);

FILL FILL_1__17208_ (
);

AND2X2 _16906_ (
    .A(_4203__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_5838_)
);

FILL FILL_0__11756_ (
);

AND2X2 _11621_ (
    .A(_1632_),
    .B(_1631_),
    .Y(_1587_[22])
);

AND2X2 _11201_ (
    .A(_1412_),
    .B(_1411_),
    .Y(_1389_[11])
);

INVX1 _19378_ (
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_8273_)
);

AND2X2 _14093_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3499_)
);

DFFSR _8828_ (
    .CLK(clk_bF$buf64),
    .D(_135_[17]),
    .Q(\datapath_1.regfile_1.regOut[3] [17]),
    .R(rst_bF$buf10),
    .S(vdd)
);

BUFX2 _8408_ (
    .A(_1_[16]),
    .Y(memoryAddress[16])
);

FILL FILL_1__13548_ (
);

AOI21X1 _12826_ (
    .A(_2389_),
    .B(_2390_),
    .C(_2388_),
    .Y(_2391_)
);

OR2X2 _12406_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .B(_2048__bF$buf4),
    .Y(_2036_)
);

AND2X2 _15298_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_4255_)
);

FILL FILL122360x251940 (
);

FILL FILL_0__16794_ (
);

FILL FILL_0__16374_ (
);

FILL FILL_1__9511_ (
);

FILL FILL345040x326040 (
);

FILL FILL411920x44460 (
);

FILL FILL57000x182780 (
);

DFFSR _8581_ (
    .CLK(clk_bF$buf91),
    .D(_3_[28]),
    .Q(\datapath_1.regfile_1.regOut[1] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL_1__18166_ (
);

FILL FILL204440x44460 (
);

FILL FILL_0__17999_ (
);

OR2X2 _17864_ (
    .A(_6749_),
    .B(_6782_),
    .Y(_6783_)
);

OR2X2 _17444_ (
    .A(_6367_),
    .B(_6368_),
    .Y(_6369_)
);

FILL FILL_0__17159_ (
);

OR2X2 _17024_ (
    .A(_5952_),
    .B(_5953_),
    .Y(_5954_)
);

FILL FILL_0__18940_ (
);

FILL FILL39520x355680 (
);

OR2X2 _9786_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_689_)
);

OR2X2 _9366_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_469_)
);

FILL FILL40280x251940 (
);

FILL FILL_0__8621_ (
);

FILL FILL187720x256880 (
);

AND2X2 _18649_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_7555_)
);

AND2X2 _18229_ (
    .A(_6326__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_7142_)
);

FILL FILL_0__13499_ (
);

AND2X2 _13784_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3252_)
);

NAND2X1 _13364_ (
    .A(_2547_),
    .B(_2902_),
    .Y(_2903_)
);

FILL FILL_0__13079_ (
);

FILL FILL_0__19305_ (
);

FILL FILL_0__14440_ (
);

FILL FILL_0__14020_ (
);

FILL FILL389880x59280 (
);

CLKBUF1 CLKBUF1_insert120 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf103)
);

CLKBUF1 CLKBUF1_insert121 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf102)
);

CLKBUF1 CLKBUF1_insert122 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf101)
);

CLKBUF1 CLKBUF1_insert123 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf100)
);

FILL FILL_0__9826_ (
);

CLKBUF1 CLKBUF1_insert124 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf99)
);

FILL FILL_0__9406_ (
);

CLKBUF1 CLKBUF1_insert125 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf98)
);

CLKBUF1 CLKBUF1_insert126 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf97)
);

FILL FILL215080x153140 (
);

CLKBUF1 CLKBUF1_insert127 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf96)
);

FILL FILL492480x291460 (
);

CLKBUF1 CLKBUF1_insert128 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf95)
);

CLKBUF1 CLKBUF1_insert129 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf94)
);

FILL FILL342760x29640 (
);

DFFSR _14989_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[8]),
    .Q(\datapath_1.mux_iord.din0 [8]),
    .R(rst_bF$buf86),
    .S(vdd)
);

AND2X2 _14569_ (
    .A(_3785_),
    .B(_3784_),
    .Y(_3738_[23])
);

OR2X2 _14149_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[2]),
    .Y(_3544_)
);

FILL FILL228000x59280 (
);

AND2X2 _15930_ (
    .A(_4877_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd2 [10])
);

FILL FILL_0__15645_ (
);

OR2X2 _15510_ (
    .A(_4462_),
    .B(_4463_),
    .Y(_4464_)
);

FILL FILL_0__10780_ (
);

FILL FILL19000x29640 (
);

FILL FILL131480x182780 (
);

DFFSR _10489_ (
    .CLK(clk_bF$buf85),
    .D(_993_[1]),
    .Q(\datapath_1.regfile_1.regOut[16] [1]),
    .R(rst_bF$buf109),
    .S(vdd)
);

OR2X2 _10069_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .B(_860__bF$buf2),
    .Y(_838_)
);

FILL FILL_1__12152_ (
);

AND2X2 _16715_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_5650_)
);

FILL FILL_0__11985_ (
);

FILL FILL171760x19760 (
);

FILL FILL_0__11565_ (
);

OR2X2 _11850_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_1745_)
);

FILL FILL50920x306280 (
);

OR2X2 _11430_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_1525_)
);

DFFSR _11010_ (
    .CLK(clk_bF$buf70),
    .D(_1257_[6]),
    .Q(\datapath_1.regfile_1.regOut[20] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

AND2X2 _19187_ (
    .A(_6317__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_8085_)
);

FILL FILL310080x370500 (
);

FILL FILL37240x217360 (
);

OR2X2 _8637_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_103_)
);

FILL FILL367840x163020 (
);

FILL FILL54720x227240 (
);

FILL FILL377720x301340 (
);

AND2X2 _12635_ (
    .A(_2199_),
    .B(_2195_),
    .Y(_2200_)
);

AND2X2 _12215_ (
    .A(_1928_),
    .B(_1927_),
    .Y(_1917_[5])
);

FILL FILL272840x123500 (
);

FILL FILL_0__13711_ (
);

FILL FILL183920x286520 (
);

BUFX2 _8390_ (
    .A(gnd),
    .Y(MemRead)
);

FILL FILL_0__14916_ (
);

FILL FILL_1__18395_ (
);

FILL FILL490960x113620 (
);

FILL FILL270560x197600 (
);

FILL FILL_0__17388_ (
);

OR2X2 _17673_ (
    .A(_6593_),
    .B(_6592_),
    .Y(_6594_)
);

AND2X2 _17253_ (
    .A(_4154__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_6180_)
);

FILL FILL126160x83980 (
);

FILL FILL115520x247000 (
);

FILL FILL414200x39520 (
);

FILL FILL_1__16708_ (
);

DFFSR _9595_ (
    .CLK(clk_bF$buf108),
    .D(_531_[10]),
    .Q(\datapath_1.regfile_1.regOut[9] [10]),
    .R(rst_bF$buf56),
    .S(vdd)
);

OR2X2 _9175_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .B(_398__bF$buf4),
    .Y(_382_)
);

FILL FILL_1__11843_ (
);

FILL FILL_0__8430_ (
);

FILL FILL_0__10836_ (
);

OR2X2 _10701_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_1159_)
);

AND2X2 _18878_ (
    .A(_6302__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_7781_)
);

FILL FILL_0_BUFX2_insert950 (
);

AND2X2 _18458_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_7367_)
);

FILL FILL_0_BUFX2_insert952 (
);

OR2X2 _18038_ (
    .A(_6953_),
    .B(_6952_),
    .Y(_6954_)
);

FILL FILL_0_BUFX2_insert953 (
);

FILL FILL_0_BUFX2_insert954 (
);

FILL FILL_0_BUFX2_insert955 (
);

AND2X2 _13593_ (
    .A(_3087__bF$buf2),
    .B(\datapath_1.ALUResult [0]),
    .Y(_3088_)
);

AND2X2 _13173_ (
    .A(_2719_),
    .B(_2722_),
    .Y(_2723_)
);

FILL FILL_0_BUFX2_insert956 (
);

FILL FILL_0_BUFX2_insert958 (
);

FILL FILL_0__19114_ (
);

FILL FILL474240x59280 (
);

FILL FILL_1__12208_ (
);

FILL FILL342000x360620 (
);

FILL FILL_0__9635_ (
);

AND2X2 _11906_ (
    .A(_1782_),
    .B(_1781_),
    .Y(_1719_[31])
);

FILL FILL133760x49400 (
);

OR2X2 _14798_ (
    .A(vdd),
    .B(_2_[14]),
    .Y(_3898_)
);

OR2X2 _14378_ (
    .A(vdd),
    .B(\datapath_1.Data [3]),
    .Y(_3678_)
);

FILL FILL_1__16461_ (
);

FILL FILL271320x4940 (
);

FILL FILL_0__15034_ (
);

AND2X2 _10298_ (
    .A(_950_),
    .B(_949_),
    .Y(_927_[11])
);

FILL FILL290320x4940 (
);

FILL FILL184680x83980 (
);

FILL FILL_0__16659_ (
);

AND2X2 _16944_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_5876_)
);

OR2X2 _16524_ (
    .A(_5460_),
    .B(_5461_),
    .Y(_5462_)
);

FILL FILL_0__16239_ (
);

OR2X2 _16104_ (
    .A(_5041_),
    .B(_5048_),
    .Y(_5049_)
);

FILL FILL_0__11374_ (
);

FILL FILL_0__17600_ (
);

FILL FILL76760x291460 (
);

FILL FILL367840x256880 (
);

OR2X2 _8866_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .B(_266__bF$buf3),
    .Y(_216_)
);

BUFX2 _8446_ (
    .A(_2_[22]),
    .Y(memoryWriteData[22])
);

FILL FILL299440x138320 (
);

OR2X2 _17729_ (
    .A(_6648_),
    .B(_6649_),
    .Y(_6650_)
);

FILL FILL454480x167960 (
);

AND2X2 _17309_ (
    .A(_6209_),
    .B(_6226_),
    .Y(_6235_)
);

FILL FILL_0__12999_ (
);

OR2X2 _12864_ (
    .A(_2422_),
    .B(_2428_),
    .Y(_2429_)
);

DFFSR _12444_ (
    .CLK(clk_bF$buf1),
    .D(_1983_[21]),
    .Q(\datapath_1.regfile_1.regOut[31] [21]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_0__12159_ (
);

OR2X2 _12024_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_1841_)
);

FILL FILL188480x0 (
);

FILL FILL_0__18805_ (
);

FILL FILL_0__13940_ (
);

FILL FILL_0__13520_ (
);

FILL FILL222680x98800 (
);

FILL FILL458280x9880 (
);

FILL FILL456760x24700 (
);

FILL FILL_0__8906_ (
);

FILL FILL188480x83980 (
);

FILL FILL156560x153140 (
);

OR2X2 _13649_ (
    .A(_3134_),
    .B(_3135_),
    .Y(_3136_)
);

OR2X2 _13229_ (
    .A(_2157__bF$buf3),
    .B(_2775_),
    .Y(_2776_)
);

FILL FILL_1__15312_ (
);

FILL FILL_0__14305_ (
);

OR2X2 _17482_ (
    .A(_6402_),
    .B(_6405_),
    .Y(_6406_)
);

OR2X2 _17062_ (
    .A(_5990_),
    .B(_5991_),
    .Y(_5992_)
);

FILL FILL25840x128440 (
);

FILL FILL433960x98800 (
);

FILL FILL_1__16937_ (
);

FILL FILL_0_CLKBUF1_insert180 (
);

FILL FILL_1__11232_ (
);

FILL FILL_0_CLKBUF1_insert181 (
);

FILL FILL_0_CLKBUF1_insert182 (
);

FILL FILL_0_CLKBUF1_insert183 (
);

FILL FILL_0_CLKBUF1_insert184 (
);

FILL FILL_0_CLKBUF1_insert186 (
);

FILL FILL265240x0 (
);

OR2X2 _10930_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_1322__bF$buf4),
    .Y(_1272_)
);

DFFSR _10510_ (
    .CLK(clk_bF$buf26),
    .D(_993_[22]),
    .Q(\datapath_1.regfile_1.regOut[16] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL_0_CLKBUF1_insert188 (
);

AND2X2 _18687_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_7593_)
);

AND2X2 _18267_ (
    .A(_6297__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_7179_)
);

FILL FILL209000x153140 (
);

FILL FILL486400x291460 (
);

FILL FILL_0__9444_ (
);

FILL FILL91960x163020 (
);

OR2X2 _11715_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_1675_)
);

FILL FILL_0__9024_ (
);

FILL FILL262960x88920 (
);

AND2X2 _14187_ (
    .A(_3569_),
    .B(_3568_),
    .Y(\datapath_1.mux_wd3.dout [14])
);

FILL FILL_0__15683_ (
);

FILL FILL_0__15263_ (
);

FILL FILL_1__8400_ (
);

FILL FILL129200x74100 (
);

FILL FILL_0__16888_ (
);

AND2X2 _16753_ (
    .A(_4236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_5688_)
);

FILL FILL_0__16468_ (
);

AND2X2 _16333_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_5274_)
);

FILL FILL409640x316160 (
);

FILL FILL_0__11183_ (
);

AND2X2 _8675_ (
    .A(_128_),
    .B(_127_),
    .Y(_69_[29])
);

FILL FILL_1__10923_ (
);

FILL FILL243200x266760 (
);

FILL FILL327560x222300 (
);

FILL FILL182400x14820 (
);

OR2X2 _17958_ (
    .A(_6867_),
    .B(_6874_),
    .Y(_6875_)
);

OR2X2 _17538_ (
    .A(_6430_),
    .B(_6461_),
    .Y(_6462_)
);

AND2X2 _17118_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_6047_)
);

OR2X2 _12673_ (
    .A(_2235_),
    .B(_2237_),
    .Y(_2238_)
);

OR2X2 _12253_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_1982__bF$buf0),
    .Y(_1954_)
);

FILL FILL338960x291460 (
);

FILL FILL_0__8715_ (
);

AND2X2 _13878_ (
    .A(_3318_),
    .B(_3317_),
    .Y(\datapath_1.alu_1.ALUInA [20])
);

AND2X2 _13458_ (
    .A(_2990_),
    .B(_2847_),
    .Y(_2991_)
);

XOR2X1 _13038_ (
    .A(_2477_),
    .B(_2475_),
    .Y(_2596_)
);

FILL FILL_1__15961_ (
);

FILL FILL_1__15541_ (
);

FILL FILL_0__14954_ (
);

FILL FILL_0__14114_ (
);

AND2X2 _17291_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_6217_)
);

FILL FILL224200x212420 (
);

FILL FILL_0__15739_ (
);

AND2X2 _15604_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_4557_)
);

FILL FILL_0__10874_ (
);

FILL FILL_0__10454_ (
);

FILL FILL361760x335920 (
);

FILL FILL235600x281580 (
);

FILL FILL250040x153140 (
);

OR2X2 _18496_ (
    .A(_7397_),
    .B(_7404_),
    .Y(_7405_)
);

OR2X2 _18076_ (
    .A(_6990_),
    .B(_6983_),
    .Y(_6991_)
);

FILL FILL_0__19152_ (
);

FILL FILL_1__12666_ (
);

AND2X2 _16809_ (
    .A(_4223__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_5743_)
);

FILL FILL232560x326040 (
);

FILL FILL_0__9673_ (
);

OR2X2 _11944_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .B(_1850__bF$buf1),
    .Y(_1788_)
);

FILL FILL_0__9253_ (
);

DFFSR _11524_ (
    .CLK(clk_bF$buf79),
    .D(_1521_[4]),
    .Q(\datapath_1.regfile_1.regOut[24] [4]),
    .R(rst_bF$buf57),
    .S(vdd)
);

OR2X2 _11104_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .B(_1388__bF$buf0),
    .Y(_1368_)
);

FILL FILL_0__12600_ (
);

FILL FILL_0__15492_ (
);

FILL FILL_0__15072_ (
);

AND2X2 _12729_ (
    .A(_2293_),
    .B(_2291_),
    .Y(_2294_)
);

DFFSR _12309_ (
    .CLK(clk_bF$buf48),
    .D(_1917_[15]),
    .Q(\datapath_1.regfile_1.regOut[30] [15]),
    .R(rst_bF$buf107),
    .S(vdd)
);

FILL FILL_0__13805_ (
);

FILL FILL_1__17284_ (
);

FILL FILL53200x375440 (
);

OR2X2 _16982_ (
    .A(_5912_),
    .B(_5911_),
    .Y(_5913_)
);

OR2X2 _16562_ (
    .A(_5498_),
    .B(_5499_),
    .Y(_5500_)
);

AND2X2 _16142_ (
    .A(_4225__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_5086_)
);

FILL FILL_1__9834_ (
);

FILL FILL298680x133380 (
);

FILL FILL234080x34580 (
);

OR2X2 _8484_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_21_)
);

FILL FILL_1__10732_ (
);

AND2X2 _17767_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_6687_)
);

OR2X2 _17347_ (
    .A(_6244__bF$buf1),
    .B(_6259__bF$buf4),
    .Y(_6273_)
);

AND2X2 _12482_ (
    .A(_2073_),
    .B(_2051_),
    .Y(_2074_)
);

DFFSR _12062_ (
    .CLK(clk_bF$buf86),
    .D(_1785_[26]),
    .Q(\datapath_1.regfile_1.regOut[28] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

FILL FILL471960x247000 (
);

FILL FILL477280x321100 (
);

FILL FILL_0__18843_ (
);

FILL FILL_0__18423_ (
);

FILL FILL_0__18003_ (
);

AND2X2 _9689_ (
    .A(_644_),
    .B(_643_),
    .Y(_597_[23])
);

AND2X2 _9269_ (
    .A(_424_),
    .B(_423_),
    .Y(_399_[12])
);

FILL FILL468920x34580 (
);

FILL FILL_0__8524_ (
);

OR2X2 _13687_ (
    .A(_3168_),
    .B(_3167_),
    .Y(_3169_)
);

NOR2X1 _13267_ (
    .A(_2800_),
    .B(_2498_),
    .Y(_2811_)
);

FILL FILL180880x59280 (
);

FILL FILL_0__14763_ (
);

FILL FILL355680x0 (
);

FILL FILL3800x242060 (
);

FILL FILL503880x301340 (
);

FILL FILL432440x291460 (
);

FILL FILL_1__11690_ (
);

OR2X2 _15833_ (
    .A(_4766_),
    .B(_4781_),
    .Y(_4782_)
);

FILL FILL_0__15548_ (
);

FILL FILL_0__15128_ (
);

OR2X2 _15413_ (
    .A(_4368_),
    .B(_4367_),
    .Y(_4369_)
);

FILL FILL_0__10683_ (
);

FILL FILL_0__10263_ (
);

FILL FILL101080x39520 (
);

FILL FILL_0__19381_ (
);

FILL FILL391400x321100 (
);

FILL FILL245480x365560 (
);

AND2X2 _16618_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_5555_)
);

FILL FILL_0__11888_ (
);

FILL FILL_1__18701_ (
);

AND2X2 _11753_ (
    .A(_1700_),
    .B(_1699_),
    .Y(_1653_[23])
);

AND2X2 _11333_ (
    .A(_1480_),
    .B(_1479_),
    .Y(_1455_[12])
);

FILL FILL432440x0 (
);

FILL FILL469680x202540 (
);

OR2X2 _9901_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_794__bF$buf1),
    .Y(_746_)
);

FILL FILL206720x182780 (
);

OR2X2 _12958_ (
    .A(_2360_),
    .B(_2350_),
    .Y(_2521_)
);

OR2X2 _12538_ (
    .A(_2127_),
    .B(_2116_),
    .Y(\control_1.next [0])
);

FILL FILL_1_BUFX2_insert884 (
);

OR2X2 _12118_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .B(_1916__bF$buf1),
    .Y(_1884_)
);

FILL FILL85120x256880 (
);

FILL FILL_1_BUFX2_insert886 (
);

FILL FILL_1_BUFX2_insert888 (
);

FILL FILL_1__14201_ (
);

FILL FILL399760x207480 (
);

FILL FILL266760x296400 (
);

OR2X2 _16791_ (
    .A(_5721_),
    .B(_5724_),
    .Y(_5725_)
);

FILL FILL232560x54340 (
);

FILL FILL_0__16086_ (
);

AND2X2 _16371_ (
    .A(_4183__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_5312_)
);

FILL FILL480320x0 (
);

FILL FILL_1__9643_ (
);

FILL FILL_1__15826_ (
);

FILL FILL_1__15406_ (
);

FILL FILL424080x14820 (
);

FILL FILL_1__10541_ (
);

FILL FILL_0__14819_ (
);

FILL FILL347320x163020 (
);

BUFX2 BUFX2_insert550 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf89)
);

BUFX2 BUFX2_insert551 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf88)
);

BUFX2 BUFX2_insert552 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf87)
);

BUFX2 BUFX2_insert553 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf86)
);

BUFX2 BUFX2_insert554 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf85)
);

AND2X2 _17996_ (
    .A(_6206__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_6912_)
);

OR2X2 _17576_ (
    .A(_6498_),
    .B(_6497_),
    .Y(_6499_)
);

BUFX2 BUFX2_insert555 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf84)
);

BUFX2 BUFX2_insert556 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf83)
);

OR2X2 _17156_ (
    .A(_6083_),
    .B(_6082_),
    .Y(_6084_)
);

BUFX2 BUFX2_insert557 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf82)
);

BUFX2 BUFX2_insert558 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf81)
);

BUFX2 BUFX2_insert559 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf80)
);

OR2X2 _12291_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_1979_)
);

FILL FILL156560x316160 (
);

FILL FILL_0__18652_ (
);

FILL FILL_0__18232_ (
);

OR2X2 _9498_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_537_)
);

DFFSR _9078_ (
    .CLK(clk_bF$buf89),
    .D(_267_[9]),
    .Q(\datapath_1.regfile_1.regOut[5] [9]),
    .R(rst_bF$buf24),
    .S(vdd)
);

FILL FILL_0__10739_ (
);

AND2X2 _10604_ (
    .A(_1114_),
    .B(_1113_),
    .Y(_1059_[27])
);

FILL FILL_0_BUFX2_insert70 (
);

FILL FILL_0_BUFX2_insert71 (
);

FILL FILL_0_BUFX2_insert72 (
);

FILL FILL_0_BUFX2_insert73 (
);

FILL FILL_0_BUFX2_insert74 (
);

FILL FILL163400x286520 (
);

FILL FILL_0_BUFX2_insert76 (
);

OR2X2 _13496_ (
    .A(ALUOut[2]),
    .B(_3079__bF$buf4),
    .Y(_3019_)
);

NAND2X1 _13076_ (
    .A(_2547_),
    .B(_2631_),
    .Y(_2632_)
);

FILL FILL_0_BUFX2_insert78 (
);

FILL FILL_0__19017_ (
);

OR2X2 _19302_ (
    .A(_8197_),
    .B(_8196_),
    .Y(_8198_)
);

FILL FILL47120x360620 (
);

FILL FILL_0__14152_ (
);

FILL FILL383040x108680 (
);

FILL FILL470440x113620 (
);

FILL FILL_0__9958_ (
);

FILL FILL_0__9538_ (
);

DFFSR _11809_ (
    .CLK(clk_bF$buf46),
    .D(_1653_[31]),
    .Q(\datapath_1.regfile_1.regOut[26] [31]),
    .R(rst_bF$buf97),
    .S(vdd)
);

FILL FILL364040x266760 (
);

FILL FILL_0__15777_ (
);

FILL FILL_0__15357_ (
);

AND2X2 _15642_ (
    .A(_4214__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_4594_)
);

OR2X2 _15222_ (
    .A(_4174_),
    .B(_4179_),
    .Y(_4180_)
);

FILL FILL_0__10072_ (
);

FILL FILL83600x29640 (
);

FILL FILL314640x4940 (
);

FILL FILL81320x286520 (
);

FILL FILL_1__17149_ (
);

FILL FILL_1__12284_ (
);

OR2X2 _16847_ (
    .A(_5779_),
    .B(_5778_),
    .Y(_5780_)
);

OR2X2 _16427_ (
    .A(_5366_),
    .B(_5365_),
    .Y(_5367_)
);

OR2X2 _16007_ (
    .A(_4952_),
    .B(_4951_),
    .Y(_4953_)
);

FILL FILL264480x345800 (
);

OR2X2 _11982_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_1813_)
);

FILL FILL_0__11697_ (
);

OR2X2 _11562_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_1593_)
);

DFFSR _11142_ (
    .CLK(clk_bF$buf24),
    .D(_1323_[9]),
    .Q(\datapath_1.regfile_1.regOut[21] [9]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_0__17923_ (
);

FILL FILL427120x306280 (
);

OR2X2 _8769_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_171_)
);

FILL FILL333640x4940 (
);

AND2X2 _9710_ (
    .A(_658_),
    .B(_657_),
    .Y(_597_[30])
);

FILL FILL_1__13489_ (
);

FILL FILL345040x212420 (
);

FILL FILL85880x24700 (
);

INVX1 _12767_ (
    .A(\datapath_1.alu_1.ALUInA [24]),
    .Y(_2332_)
);

AND2X2 _12347_ (
    .A(_1996_),
    .B(_1995_),
    .Y(_1983_[6])
);

FILL FILL430920x340860 (
);

FILL FILL_0__18708_ (
);

FILL FILL_0__13423_ (
);

FILL FILL_0__13003_ (
);

FILL FILL352640x4940 (
);

AND2X2 _16180_ (
    .A(_4241__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_5124_)
);

FILL FILL291080x69160 (
);

FILL FILL_0__8809_ (
);

FILL FILL193040x123500 (
);

FILL FILL_0__14628_ (
);

OR2X2 _14913_ (
    .A(\datapath_1.mux_pcsrc.dout [9]),
    .B(_4001__bF$buf4),
    .Y(_3955_)
);

FILL FILL_0__14208_ (
);

NOR2X1 _17385_ (
    .A(_6310__bF$buf2),
    .B(_6307_),
    .Y(_6311_)
);

FILL FILL_0__18881_ (
);

FILL FILL256880x360620 (
);

FILL FILL_0__18041_ (
);

FILL FILL89680x24700 (
);

FILL FILL_1__11975_ (
);

FILL FILL314640x143260 (
);

FILL FILL_0__10968_ (
);

OR2X2 _10833_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_1227_)
);

FILL FILL_0__10548_ (
);

OR2X2 _10413_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_1007_)
);

DFFSR _19531_ (
    .CLK(clk_bF$buf98),
    .D(_8320_[8]),
    .Q(\datapath_1.regfile_1.regOut[0] [8]),
    .R(rst_bF$buf87),
    .S(vdd)
);

FILL FILL_0__19246_ (
);

AND2X2 _19111_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_8010_)
);

FILL FILL_0__9767_ (
);

AND2X2 _11618_ (
    .A(_1630_),
    .B(_1629_),
    .Y(_1587_[21])
);

FILL FILL130720x266760 (
);

FILL FILL50160x232180 (
);

FILL FILL136040x340860 (
);

FILL FILL117040x177840 (
);

AND2X2 _15871_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_4819_)
);

FILL FILL_0__15586_ (
);

AND2X2 _15451_ (
    .A(_4239__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_4406_)
);

NOR2X1 _15031_ (
    .A(_4019_),
    .B(\datapath_1.a3 [3]),
    .Y(_4020_)
);

FILL FILL354920x103740 (
);

FILL FILL_1__17798_ (
);

FILL FILL383800x0 (
);

FILL FILL_1__17378_ (
);

FILL FILL_1__12093_ (
);

OR2X2 _16656_ (
    .A(_5588_),
    .B(_5591_),
    .Y(_5592_)
);

AND2X2 _16236_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_5179_)
);

DFFSR _11791_ (
    .CLK(clk_bF$buf85),
    .D(_1653_[13]),
    .Q(\datapath_1.regfile_1.regOut[26] [13]),
    .R(rst_bF$buf109),
    .S(vdd)
);

OR2X2 _11371_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .B(_1520__bF$buf0),
    .Y(_1506_)
);

FILL FILL_1__9928_ (
);

FILL FILL148960x148200 (
);

FILL FILL170240x266760 (
);

FILL FILL_0__17312_ (
);

OR2X2 _8998_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .B(_332__bF$buf1),
    .Y(_284_)
);

DFFSR _8578_ (
    .CLK(clk_bF$buf16),
    .D(_3_[25]),
    .Q(\datapath_1.regfile_1.regOut[1] [25]),
    .R(rst_bF$buf20),
    .S(vdd)
);

FILL FILL352640x177840 (
);

OR2X2 _12996_ (
    .A(_2321_),
    .B(_2556_),
    .Y(_2557_)
);

OR2X2 _12576_ (
    .A(\control_1.next [1]),
    .B(_2145_),
    .Y(_2148_)
);

OR2X2 _12156_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_1909_)
);

FILL FILL_0__18937_ (
);

OR2X2 _18802_ (
    .A(_7705_),
    .B(_7704_),
    .Y(_7706_)
);

FILL FILL_0__18517_ (
);

FILL FILL_0__13652_ (
);

FILL FILL_0__13232_ (
);

FILL FILL52440x187720 (
);

FILL FILL_0__8618_ (
);

FILL FILL_1__9261_ (
);

BUFX2 BUFX2_insert1110 (
    .A(_1454_),
    .Y(_1454__bF$buf4)
);

BUFX2 BUFX2_insert1111 (
    .A(_1454_),
    .Y(_1454__bF$buf3)
);

BUFX2 BUFX2_insert1112 (
    .A(_1454_),
    .Y(_1454__bF$buf2)
);

BUFX2 BUFX2_insert1113 (
    .A(_1454_),
    .Y(_1454__bF$buf1)
);

BUFX2 BUFX2_insert1114 (
    .A(_1454_),
    .Y(_1454__bF$buf0)
);

FILL FILL462080x172900 (
);

BUFX2 BUFX2_insert1115 (
    .A(_2048_),
    .Y(_2048__bF$buf4)
);

BUFX2 BUFX2_insert1116 (
    .A(_2048_),
    .Y(_2048__bF$buf3)
);

BUFX2 BUFX2_insert1117 (
    .A(_2048_),
    .Y(_2048__bF$buf2)
);

FILL FILL66880x148200 (
);

BUFX2 BUFX2_insert1118 (
    .A(_2048_),
    .Y(_2048__bF$buf1)
);

BUFX2 BUFX2_insert1119 (
    .A(_2048_),
    .Y(_2048__bF$buf0)
);

AND2X2 _14722_ (
    .A(_3867_),
    .B(_3866_),
    .Y(_3804_[31])
);

AND2X2 _14302_ (
    .A(_3647_),
    .B(_3646_),
    .Y(_3606_[20])
);

BUFX2 BUFX2_insert930 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf2 )
);

BUFX2 BUFX2_insert931 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf1 )
);

BUFX2 BUFX2_insert932 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf0 )
);

BUFX2 BUFX2_insert933 (
    .A(_3089_),
    .Y(_3089__bF$buf4)
);

BUFX2 BUFX2_insert934 (
    .A(_3089_),
    .Y(_3089__bF$buf3)
);

BUFX2 BUFX2_insert935 (
    .A(_3089_),
    .Y(_3089__bF$buf2)
);

BUFX2 BUFX2_insert936 (
    .A(_3089_),
    .Y(_3089__bF$buf1)
);

AND2X2 _17194_ (
    .A(_4146__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_6122_)
);

BUFX2 BUFX2_insert937 (
    .A(_3089_),
    .Y(_3089__bF$buf0)
);

FILL FILL415720x217360 (
);

BUFX2 BUFX2_insert938 (
    .A(_6287_),
    .Y(_6287__bF$buf4)
);

BUFX2 BUFX2_insert939 (
    .A(_6287_),
    .Y(_6287__bF$buf3)
);

FILL FILL_0__18270_ (
);

FILL FILL_1__16229_ (
);

FILL FILL438520x301340 (
);

OR2X2 _15927_ (
    .A(_4874_),
    .B(_4867_),
    .Y(_4875_)
);

OR2X2 _15507_ (
    .A(_4459_),
    .B(_4460_),
    .Y(_4461_)
);

DFFSR _10642_ (
    .CLK(clk_bF$buf81),
    .D(_1059_[25]),
    .Q(\datapath_1.regfile_1.regOut[17] [25]),
    .R(rst_bF$buf13),
    .S(vdd)
);

OR2X2 _10222_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .B(_926__bF$buf0),
    .Y(_920_)
);

FILL FILL419520x138320 (
);

OR2X2 _18399_ (
    .A(_7305_),
    .B(_7308_),
    .Y(_7309_)
);

FILL FILL368600x306280 (
);

OR2X2 _19340_ (
    .A(_8235_),
    .B(_8232_),
    .Y(_8236_)
);

FILL FILL_1__12989_ (
);

FILL FILL_0__9576_ (
);

FILL FILL_0__9156_ (
);

OR2X2 _11847_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .Y(_1743_)
);

OR2X2 _11427_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_1523_)
);

DFFSR _11007_ (
    .CLK(clk_bF$buf57),
    .D(_1257_[3]),
    .Q(\datapath_1.regfile_1.regOut[20] [3]),
    .R(rst_bF$buf81),
    .S(vdd)
);

FILL FILL_1__13930_ (
);

FILL FILL111720x69160 (
);

FILL FILL_0__12923_ (
);

FILL FILL481080x158080 (
);

FILL FILL_0__12503_ (
);

FILL FILL297920x281580 (
);

OR2X2 _15680_ (
    .A(_4630_),
    .B(_4629_),
    .Y(_4631_)
);

FILL FILL280440x365560 (
);

FILL FILL373160x123500 (
);

AND2X2 _15260_ (
    .A(_4217__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_4218_)
);

FILL FILL_1__8532_ (
);

FILL FILL303240x29640 (
);

OR2X2 _16885_ (
    .A(_5817_),
    .B(_5816_),
    .Y(_5818_)
);

AND2X2 _16465_ (
    .A(_4214__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_5404_)
);

AND2X2 _16045_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_4991_)
);

AND2X2 _11180_ (
    .A(_1398_),
    .B(_1397_),
    .Y(_1389_[4])
);

FILL FILL_0__17961_ (
);

FILL FILL_0__17541_ (
);

FILL FILL_0__17121_ (
);

FILL FILL132240x19760 (
);

OR2X2 _12385_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .B(_2048__bF$buf0),
    .Y(_2022_)
);

FILL FILL_0__18746_ (
);

AND2X2 _18611_ (
    .A(_6282__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_7518_)
);

FILL FILL_0__13881_ (
);

FILL FILL_0__13041_ (
);

FILL FILL310840x266760 (
);

FILL FILL347320x326040 (
);

FILL FILL_0__8847_ (
);

FILL FILL_0__8427_ (
);

FILL FILL191520x316160 (
);

FILL FILL227240x44460 (
);

FILL FILL259160x291460 (
);

OR2X2 _14951_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [22]),
    .Y(_3980_)
);

FILL FILL_0__14246_ (
);

OR2X2 _14531_ (
    .A(IRWrite_bF$buf3),
    .B(\datapath_1.PCJump [13]),
    .Y(_3760_)
);

AND2X2 _14111_ (
    .A(_3352__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3515_)
);

FILL FILL18240x14820 (
);

FILL FILL_1__16878_ (
);

FILL FILL_1__11593_ (
);

OR2X2 _15736_ (
    .A(_4671_),
    .B(_4686_),
    .Y(_4687_)
);

AND2X2 _15316_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_4273_)
);

FILL FILL_0__10586_ (
);

AND2X2 _10871_ (
    .A(_1252_),
    .B(_1251_),
    .Y(_1191_[30])
);

AND2X2 _10451_ (
    .A(_1032_),
    .B(_1031_),
    .Y(_993_[19])
);

AND2X2 _10031_ (
    .A(_812_),
    .B(_811_),
    .Y(_795_[8])
);

BUFX2 BUFX2_insert80 (
    .A(_1718_),
    .Y(_1718__bF$buf4)
);

BUFX2 BUFX2_insert81 (
    .A(_1718_),
    .Y(_1718__bF$buf3)
);

BUFX2 BUFX2_insert82 (
    .A(_1718_),
    .Y(_1718__bF$buf2)
);

BUFX2 BUFX2_insert83 (
    .A(_1718_),
    .Y(_1718__bF$buf1)
);

BUFX2 BUFX2_insert84 (
    .A(_1718_),
    .Y(_1718__bF$buf0)
);

FILL FILL_0__16812_ (
);

BUFX2 BUFX2_insert85 (
    .A(_3079_),
    .Y(_3079__bF$buf4)
);

BUFX2 BUFX2_insert86 (
    .A(_3079_),
    .Y(_3079__bF$buf3)
);

BUFX2 BUFX2_insert87 (
    .A(_3079_),
    .Y(_3079__bF$buf2)
);

FILL FILL468920x350740 (
);

BUFX2 BUFX2_insert88 (
    .A(_3079_),
    .Y(_3079__bF$buf1)
);

FILL FILL483360x222300 (
);

BUFX2 BUFX2_insert89 (
    .A(_3079_),
    .Y(_3079__bF$buf0)
);

FILL FILL_0__19284_ (
);

FILL FILL_0__9385_ (
);

DFFSR _11656_ (
    .CLK(clk_bF$buf66),
    .D(_1587_[7]),
    .Q(\datapath_1.regfile_1.regOut[25] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

OR2X2 _11236_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .B(_1454__bF$buf0),
    .Y(_1436_)
);

FILL FILL147440x158080 (
);

FILL FILL158080x29640 (
);

OR2X2 _9804_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_701_)
);

FILL FILL_0__13937_ (
);

FILL FILL_0__13517_ (
);

AND2X2 _13802_ (
    .A(_3084__bF$buf3),
    .B(\datapath_1.PCJump [30]),
    .Y(_3267_)
);

OR2X2 _16694_ (
    .A(_5626_),
    .B(_5629_),
    .Y(_5630_)
);

FILL FILL312360x370500 (
);

FILL FILL340480x103740 (
);

FILL FILL36480x64220 (
);

AND2X2 _16274_ (
    .A(_4172__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_5216_)
);

FILL FILL39520x217360 (
);

FILL FILL426360x118560 (
);

FILL FILL_1__9546_ (
);

FILL FILL_0__17770_ (
);

FILL FILL_0__17350_ (
);

FILL FILL391400x281580 (
);

FILL FILL_1__10864_ (
);

OR2X2 _17899_ (
    .A(_6815_),
    .B(_6816_),
    .Y(_6817_)
);

AND2X2 _17479_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_6403_)
);

FILL FILL21280x271700 (
);

OR2X2 _17059_ (
    .A(_5988_),
    .B(_5987_),
    .Y(_5989_)
);

FILL FILL_1__19142_ (
);

DFFSR _12194_ (
    .CLK(clk_bF$buf11),
    .D(_1851_[29]),
    .Q(\datapath_1.regfile_1.regOut[29] [29]),
    .R(rst_bF$buf111),
    .S(vdd)
);

AND2X2 _18840_ (
    .A(_7743_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.rd1 [22])
);

FILL FILL_0__18135_ (
);

AND2X2 _18420_ (
    .A(_6262__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_7330_)
);

FILL FILL443080x355680 (
);

AND2X2 _18000_ (
    .A(_6221__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_6916_)
);

FILL FILL_0__13690_ (
);

FILL FILL_0__13270_ (
);

FILL FILL_0__8656_ (
);

FILL FILL255360x187720 (
);

OR2X2 _10927_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .B(_1322__bF$buf4),
    .Y(_1270_)
);

DFFSR _10507_ (
    .CLK(clk_bF$buf86),
    .D(_993_[19]),
    .Q(\datapath_1.regfile_1.regOut[16] [19]),
    .R(rst_bF$buf72),
    .S(vdd)
);

INVX1 _13399_ (
    .A(_2935_),
    .Y(\datapath_1.ALUResult [3])
);

FILL FILL505400x153140 (
);

FILL FILL417240x24700 (
);

OR2X2 _19205_ (
    .A(_8101_),
    .B(_8102_),
    .Y(_8103_)
);

FILL FILL272840x197600 (
);

OR2X2 _14760_ (
    .A(\datapath_1.rd2 [1]),
    .B(_3935__bF$buf3),
    .Y(_3873_)
);

DFFSR _14340_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[4]),
    .Q(ALUOut[4]),
    .R(rst_bF$buf29),
    .S(vdd)
);

FILL FILL117800x247000 (
);

FILL FILL421800x182780 (
);

FILL FILL57760x88920 (
);

FILL FILL_1__16267_ (
);

AND2X2 _15965_ (
    .A(_4241__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_4912_)
);

OR2X2 _15545_ (
    .A(_4467_),
    .B(_4498_),
    .Y(_4499_)
);

NAND3X1 _15125_ (
    .A(_4031_),
    .B(_4002_),
    .C(_4017_),
    .Y(_4102_)
);

FILL FILL_0__10395_ (
);

OR2X2 _10680_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_1145_)
);

DFFSR _10260_ (
    .CLK(clk_bF$buf108),
    .D(_861_[30]),
    .Q(\datapath_1.regfile_1.regOut[14] [30]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL_0__16621_ (
);

FILL FILL243960x281580 (
);

FILL FILL_0__19093_ (
);

FILL FILL266000x29640 (
);

FILL FILL354160x306280 (
);

FILL FILL441560x311220 (
);

AND2X2 _11885_ (
    .A(_1768_),
    .B(_1767_),
    .Y(_1719_[24])
);

AND2X2 _11465_ (
    .A(_1548_),
    .B(_1547_),
    .Y(_1521_[13])
);

AND2X2 _11045_ (
    .A(_1328_),
    .B(_1327_),
    .Y(_1323_[2])
);

FILL FILL_0__17826_ (
);

FILL FILL35720x247000 (
);

FILL FILL_0__17406_ (
);

FILL FILL_0__12121_ (
);

FILL FILL370120x44460 (
);

DFFSR _9613_ (
    .CLK(clk_bF$buf91),
    .D(_531_[28]),
    .Q(\datapath_1.regfile_1.regOut[9] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL253080x370500 (
);

FILL FILL268280x24700 (
);

FILL FILL_0__13746_ (
);

FILL FILL_0__13326_ (
);

OR2X2 _13611_ (
    .A(_3103_),
    .B(_3100_),
    .Y(\datapath_1.mux_pcsrc.dout [2])
);

OR2X2 _16083_ (
    .A(_5026_),
    .B(_5027_),
    .Y(_5028_)
);

FILL FILL6080x138320 (
);

FILL FILL_1__10673_ (
);

OR2X2 _14816_ (
    .A(vdd),
    .B(_2_[20]),
    .Y(_3910_)
);

AND2X2 _17288_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_6214_)
);

FILL FILL_0__18784_ (
);

FILL FILL_0__18364_ (
);

FILL FILL_1__11878_ (
);

FILL FILL_1__11038_ (
);

FILL FILL379240x345800 (
);

FILL FILL_0__8465_ (
);

AND2X2 _10736_ (
    .A(_1182_),
    .B(_1181_),
    .Y(_1125_[28])
);

AND2X2 _10316_ (
    .A(_962_),
    .B(_961_),
    .Y(_927_[17])
);

FILL FILL_0__11812_ (
);

OR2X2 _19434_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8325_)
);

FILL FILL_0__19149_ (
);

OR2X2 _19014_ (
    .A(_7911_),
    .B(_7914_),
    .Y(_7915_)
);

FILL FILL_1__16496_ (
);

FILL FILL102600x59280 (
);

AND2X2 _15774_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_4724_)
);

FILL FILL_0__15489_ (
);

AND2X2 _15354_ (
    .A(_4310_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.rd2 [1])
);

FILL FILL_0__15069_ (
);

FILL FILL_1__8626_ (
);

FILL FILL_0__16430_ (
);

FILL FILL44840x365560 (
);

FILL FILL_0__16010_ (
);

OR2X2 _16979_ (
    .A(_5909_),
    .B(_5908_),
    .Y(_5910_)
);

OR2X2 _16559_ (
    .A(_5496_),
    .B(_5493_),
    .Y(_5497_)
);

AND2X2 _16139_ (
    .A(_4130__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_5083_)
);

OR2X2 _11694_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_1661_)
);

FILL FILL_1__18642_ (
);

DFFSR _11274_ (
    .CLK(clk_bF$buf113),
    .D(_1389_[12]),
    .Q(\datapath_1.regfile_1.regOut[22] [12]),
    .R(rst_bF$buf102),
    .S(vdd)
);

FILL FILL435480x187720 (
);

AND2X2 _17920_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_6838_)
);

FILL FILL_0__17635_ (
);

FILL FILL_0__17215_ (
);

AND2X2 _17500_ (
    .A(_6321__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_6424_)
);

FILL FILL_0__12770_ (
);

FILL FILL_1__10309_ (
);

AND2X2 _9842_ (
    .A(_726_),
    .B(_725_),
    .Y(_663_[31])
);

AND2X2 _9422_ (
    .A(_506_),
    .B(_505_),
    .Y(_465_[20])
);

AND2X2 _9002_ (
    .A(_286_),
    .B(_285_),
    .Y(_267_[9])
);

FILL FILL205960x291460 (
);

FILL FILL505400x19760 (
);

AND2X2 _12899_ (
    .A(_2461_),
    .B(_2463_),
    .Y(_2464_)
);

OR2X2 _12479_ (
    .A(_2071_),
    .B(_2066_),
    .Y(ALUControl[1])
);

FILL FILL_1__19427_ (
);

DFFSR _12059_ (
    .CLK(clk_bF$buf101),
    .D(_1785_[23]),
    .Q(\datapath_1.regfile_1.regOut[28] [23]),
    .R(rst_bF$buf89),
    .S(vdd)
);

FILL FILL_1__19007_ (
);

OR2X2 _18705_ (
    .A(_7607_),
    .B(_7610_),
    .Y(_7611_)
);

FILL FILL_0__13975_ (
);

OR2X2 _13840_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [8]),
    .Y(_3293_)
);

FILL FILL_0__13555_ (
);

AND2X2 _13420_ (
    .A(_2954_),
    .B(_2953_),
    .Y(_2955_)
);

AND2X2 _13000_ (
    .A(_2560_),
    .B(_2546_),
    .Y(_2561_)
);

FILL FILL_1__15347_ (
);

FILL FILL_1__10062_ (
);

FILL FILL108680x54340 (
);

DFFSR _14625_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[31]),
    .Q(\control_1.op [5]),
    .R(rst_bF$buf100),
    .S(vdd)
);

AND2X2 _14205_ (
    .A(_3581_),
    .B(_3580_),
    .Y(\datapath_1.mux_wd3.dout [20])
);

OR2X2 _17097_ (
    .A(_6018_),
    .B(_6025_),
    .Y(_6026_)
);

FILL FILL163400x172900 (
);

FILL FILL_1__19180_ (
);

FILL FILL_0__18593_ (
);

FILL FILL260680x123500 (
);

FILL FILL154280x276640 (
);

OR2X2 _10965_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_1295_)
);

OR2X2 _10545_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_1075_)
);

DFFSR _10125_ (
    .CLK(clk_bF$buf8),
    .D(_795_[24]),
    .Q(\datapath_1.regfile_1.regOut[13] [24]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL_0__16906_ (
);

FILL FILL_0__11201_ (
);

FILL FILL_0__19378_ (
);

FILL FILL171760x286520 (
);

FILL FILL319960x54340 (
);

OR2X2 _19243_ (
    .A(_8138_),
    .B(_8139_),
    .Y(_8140_)
);

FILL FILL_0__14093_ (
);

FILL FILL276640x0 (
);

FILL FILL357200x98800 (
);

FILL FILL_0__9899_ (
);

FILL FILL_0__9059_ (
);

FILL FILL_1__13413_ (
);

FILL FILL_0__12406_ (
);

FILL FILL252320x153140 (
);

FILL FILL_0__15298_ (
);

OR2X2 _15583_ (
    .A(_4534_),
    .B(_4535_),
    .Y(_4536_)
);

NAND2X1 _15163_ (
    .A(RegWrite),
    .B(_4124_),
    .Y(_4125_)
);

FILL FILL217360x316160 (
);

FILL FILL234840x326040 (
);

FILL FILL135280x222300 (
);

FILL FILL224200x286520 (
);

AND2X2 _16788_ (
    .A(_4151__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_5722_)
);

AND2X2 _16368_ (
    .A(_4217__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_5309_)
);

OR2X2 _11083_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .B(_1388__bF$buf3),
    .Y(_1354_)
);

FILL FILL_1__18031_ (
);

FILL FILL393680x197600 (
);

FILL FILL321480x237120 (
);

FILL FILL_0__17864_ (
);

FILL FILL238640x247000 (
);

FILL FILL34960x108680 (
);

OR2X2 _9651_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_619_)
);

INVX2 _9231_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .Y(_464_)
);

OR2X2 _12288_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_1977_)
);

FILL FILL63840x44460 (
);

FILL FILL_1__14791_ (
);

FILL FILL_0__18649_ (
);

OR2X2 _18934_ (
    .A(_7835_),
    .B(_7822_),
    .Y(_7836_)
);

FILL FILL_0__18229_ (
);

OR2X2 _18514_ (
    .A(_7389_),
    .B(_7422_),
    .Y(_7423_)
);

FILL FILL464360x34580 (
);

FILL FILL_0__13364_ (
);

FILL FILL216600x54340 (
);

FILL FILL_1__9393_ (
);

FILL FILL123880x24700 (
);

FILL FILL_1__15996_ (
);

DFFSR _14854_ (
    .CLK(clk_bF$buf58),
    .D(_3870_[2]),
    .Q(_2_[2]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__14569_ (
);

FILL FILL395200x365560 (
);

AND2X2 _14434_ (
    .A(_3715_),
    .B(_3714_),
    .Y(_3672_[21])
);

OR2X2 _14014_ (
    .A(_3431_),
    .B(_3430_),
    .Y(_3432_)
);

FILL FILL_0__15930_ (
);

FILL FILL104120x251940 (
);

FILL FILL_0__15510_ (
);

FILL FILL492480x316160 (
);

FILL FILL67640x44460 (
);

OR2X2 _15639_ (
    .A(_4590_),
    .B(_4587_),
    .Y(_4591_)
);

NOR3X1 _15219_ (
    .A(_4145_),
    .B(_4144_),
    .C(_4150_),
    .Y(_4177_)
);

FILL FILL468160x34580 (
);

DFFSR _10774_ (
    .CLK(clk_bF$buf110),
    .D(_1125_[28]),
    .Q(\datapath_1.regfile_1.regOut[18] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

OR2X2 _10354_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .B(_992__bF$buf3),
    .Y(_988_)
);

FILL FILL235600x330980 (
);

FILL FILL20520x14820 (
);

FILL FILL408880x158080 (
);

FILL FILL_0__11850_ (
);

FILL FILL_0__11430_ (
);

FILL FILL127680x24700 (
);

FILL FILL_0__19187_ (
);

OR2X2 _19472_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_8350_)
);

AND2X2 _19052_ (
    .A(_6247__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_7952_)
);

OR2X2 _8922_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_253_)
);

OR2X2 _8502_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_33_)
);

OR2X2 _11979_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_1811_)
);

FILL FILL_0__9288_ (
);

OR2X2 _11559_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_1591_)
);

FILL FILL_1__18507_ (
);

DFFSR _11139_ (
    .CLK(clk_bF$buf7),
    .D(_1323_[6]),
    .Q(\datapath_1.regfile_1.regOut[21] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

NAND2X1 _12920_ (
    .A(_2360_),
    .B(_2356_),
    .Y(_2485_)
);

FILL FILL_0__12635_ (
);

FILL FILL_0__12215_ (
);

NOR3X1 _12500_ (
    .A(_2097_),
    .B(\control_1.reg_state.dout [1]),
    .C(\control_1.reg_state.dout [0]),
    .Y(PCSource[1])
);

FILL FILL_1_BUFX2_insert505 (
);

FILL FILL_1_BUFX2_insert507 (
);

FILL FILL_1_BUFX2_insert509 (
);

OR2X2 _15392_ (
    .A(_4347_),
    .B(_4344_),
    .Y(_4348_)
);

AND2X2 _9707_ (
    .A(_656_),
    .B(_655_),
    .Y(_597_[29])
);

FILL FILL275120x330980 (
);

FILL FILL_1__8664_ (
);

FILL FILL266760x207480 (
);

FILL FILL_1__14427_ (
);

FILL FILL503880x375440 (
);

OR2X2 _13705_ (
    .A(_3182_),
    .B(_3183_),
    .Y(_3184_)
);

AND2X2 _16597_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [21]),
    .Y(_5534_)
);

AND2X2 _16177_ (
    .A(_4236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_5121_)
);

FILL FILL_1__18680_ (
);

FILL FILL_1__18260_ (
);

FILL FILL_0__17253_ (
);

OR2X2 _9880_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .B(_794__bF$buf2),
    .Y(_732_)
);

DFFSR _9460_ (
    .CLK(clk_bF$buf73),
    .D(_465_[4]),
    .Q(\datapath_1.regfile_1.regOut[8] [4]),
    .R(rst_bF$buf39),
    .S(vdd)
);

OR2X2 _9040_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_332__bF$buf4),
    .Y(_312_)
);

FILL FILL462840x54340 (
);

OR2X2 _12097_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .B(_1916__bF$buf3),
    .Y(_1870_)
);

FILL FILL_0__10701_ (
);

FILL FILL_0__18878_ (
);

AND2X2 _18743_ (
    .A(_6317__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_7648_)
);

FILL FILL_0__18458_ (
);

OR2X2 _18323_ (
    .A(_7233_),
    .B(_7232_),
    .Y(_7234_)
);

FILL FILL_0__13593_ (
);

FILL FILL_0__8979_ (
);

FILL FILL_1__12913_ (
);

FILL FILL349600x163020 (
);

FILL FILL_0__9920_ (
);

FILL FILL_0__11906_ (
);

FILL FILL_1__15385_ (
);

FILL FILL345800x108680 (
);

FILL FILL138320x93860 (
);

FILL FILL322240x93860 (
);

DFFSR _19528_ (
    .CLK(clk_bF$buf49),
    .D(_8320_[5]),
    .Q(\datapath_1.regfile_1.regOut[0] [5]),
    .R(rst_bF$buf106),
    .S(vdd)
);

AND2X2 _19108_ (
    .A(_6229__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_8007_)
);

FILL FILL_0__14798_ (
);

OR2X2 _14663_ (
    .A(vdd),
    .B(\datapath_1.a [12]),
    .Y(_3828_)
);

FILL FILL_0__14378_ (
);

OR2X2 _14243_ (
    .A(vdd),
    .B(ALUOut[1]),
    .Y(_3608_)
);

FILL FILL158840x316160 (
);

FILL FILL23560x98800 (
);

AND2X2 _15868_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_4816_)
);

OR2X2 _15448_ (
    .A(_4395_),
    .B(_4402_),
    .Y(_4403_)
);

INVX1 _15028_ (
    .A(\datapath_1.a3 [4]),
    .Y(_4017_)
);

AND2X2 _10583_ (
    .A(_1100_),
    .B(_1099_),
    .Y(_1059_[20])
);

AND2X2 _10163_ (
    .A(_880_),
    .B(_879_),
    .Y(_861_[9])
);

FILL FILL393680x39520 (
);

FILL FILL271320x360620 (
);

FILL FILL_0__16944_ (
);

FILL FILL_0__16104_ (
);

FILL FILL49400x360620 (
);

FILL FILL385320x108680 (
);

AND2X2 _19281_ (
    .A(_6232__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_8178_)
);

OR2X2 _8731_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .B(_200__bF$buf3),
    .Y(_146_)
);

FILL FILL366320x266760 (
);

DFFSR _11788_ (
    .CLK(clk_bF$buf76),
    .D(_1653_[10]),
    .Q(\datapath_1.regfile_1.regOut[26] [10]),
    .R(rst_bF$buf110),
    .S(vdd)
);

OR2X2 _11368_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_1520__bF$buf0),
    .Y(_1504_)
);

FILL FILL_1__13871_ (
);

FILL FILL_0__17729_ (
);

FILL FILL_0__12864_ (
);

FILL FILL_0__12024_ (
);

FILL FILL389120x350740 (
);

FILL FILL311600x316160 (
);

FILL FILL300200x0 (
);

OR2X2 _9936_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_769_)
);

FILL FILL27360x98800 (
);

OR2X2 _9516_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_549_)
);

FILL FILL_1__8473_ (
);

FILL FILL83600x286520 (
);

FILL FILL223440x281580 (
);

FILL FILL_1__14236_ (
);

OR2X2 _13934_ (
    .A(_3361_),
    .B(_3362_),
    .Y(_3363_)
);

FILL FILL266760x345800 (
);

OR2X2 _13514_ (
    .A(ALUOut[8]),
    .B(_3079__bF$buf3),
    .Y(_3031_)
);

FILL FILL123120x375440 (
);

FILL FILL_1__9678_ (
);

BUFX2 BUFX2_insert1080 (
    .A(_4200_),
    .Y(_4200__bF$buf4)
);

BUFX2 BUFX2_insert1081 (
    .A(_4200_),
    .Y(_4200__bF$buf3)
);

BUFX2 BUFX2_insert1082 (
    .A(_4200_),
    .Y(_4200__bF$buf2)
);

FILL FILL_0__17482_ (
);

BUFX2 BUFX2_insert1083 (
    .A(_4200_),
    .Y(_4200__bF$buf1)
);

BUFX2 BUFX2_insert1084 (
    .A(_4200_),
    .Y(_4200__bF$buf0)
);

BUFX2 BUFX2_insert1085 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf4 )
);

BUFX2 BUFX2_insert1086 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf3 )
);

BUFX2 BUFX2_insert1087 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf2 )
);

BUFX2 BUFX2_insert1088 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf1 )
);

BUFX2 BUFX2_insert1089 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf0 )
);

FILL FILL_1__10996_ (
);

AND2X2 _14719_ (
    .A(_3865_),
    .B(_3864_),
    .Y(_3804_[30])
);

FILL FILL347320x212420 (
);

FILL FILL_1__16802_ (
);

FILL FILL270560x24700 (
);

FILL FILL_1_CLKBUF1_insert211 (
);

FILL FILL_1_CLKBUF1_insert213 (
);

FILL FILL_1_CLKBUF1_insert215 (
);

FILL FILL_0__18687_ (
);

AND2X2 _18972_ (
    .A(_6211__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_7873_)
);

OR2X2 _18552_ (
    .A(_7459_),
    .B(_7458_),
    .Y(_7460_)
);

FILL FILL_0__18267_ (
);

FILL FILL384560x93860 (
);

OR2X2 _18132_ (
    .A(_7042_),
    .B(_7045_),
    .Y(_7046_)
);

FILL FILL_0__8788_ (
);

DFFSR _10639_ (
    .CLK(clk_bF$buf26),
    .D(_1059_[22]),
    .Q(\datapath_1.regfile_1.regOut[17] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

OR2X2 _10219_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .B(_926__bF$buf4),
    .Y(_918_)
);

FILL FILL_0__11715_ (
);

FILL FILL345040x286520 (
);

AND2X2 _19337_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_8233_)
);

OR2X2 _14892_ (
    .A(\datapath_1.mux_pcsrc.dout [2]),
    .B(_4001__bF$buf1),
    .Y(_3941_)
);

FILL FILL_0__14187_ (
);

DFFSR _14472_ (
    .CLK(clk_bF$buf78),
    .D(_3672_[7]),
    .Q(\datapath_1.Data [7]),
    .R(rst_bF$buf85),
    .S(vdd)
);

AND2X2 _14052_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3464_)
);

FILL FILL362520x296400 (
);

FILL FILL12920x232180 (
);

OR2X2 _15677_ (
    .A(_4626_),
    .B(_4627_),
    .Y(_4628_)
);

FILL FILL193040x197600 (
);

AND2X2 _15257_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_4215_)
);

FILL FILL221920x103740 (
);

FILL FILL_1__17760_ (
);

INVX2 _10392_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .Y(_1058_)
);

FILL FILL_0__16753_ (
);

FILL FILL_0__16333_ (
);

AND2X2 _19090_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_7990_)
);

FILL FILL342000x182780 (
);

DFFSR _8960_ (
    .CLK(clk_bF$buf83),
    .D(_201_[20]),
    .Q(\datapath_1.regfile_1.regOut[4] [20]),
    .R(rst_bF$buf17),
    .S(vdd)
);

AND2X2 _8540_ (
    .A(_58_),
    .B(_57_),
    .Y(_3_[27])
);

FILL FILL52440x232180 (
);

FILL FILL138320x340860 (
);

AND2X2 _11597_ (
    .A(_1616_),
    .B(_1615_),
    .Y(_1587_[14])
);

FILL FILL_1__18125_ (
);

AND2X2 _11177_ (
    .A(_1396_),
    .B(_1395_),
    .Y(_1389_[3])
);

FILL FILL_0__17958_ (
);

AND2X2 _17823_ (
    .A(_6262__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_6742_)
);

AND2X2 _17403_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_6329_)
);

FILL FILL_0__17118_ (
);

FILL FILL_0__12673_ (
);

FILL FILL_0__12253_ (
);

DFFSR _9745_ (
    .CLK(clk_bF$buf95),
    .D(_597_[31]),
    .Q(\datapath_1.regfile_1.regOut[10] [31]),
    .R(rst_bF$buf30),
    .S(vdd)
);

OR2X2 _9325_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .B(_464__bF$buf3),
    .Y(_462_)
);

OR2X2 _18608_ (
    .A(_7511_),
    .B(_7514_),
    .Y(_7515_)
);

FILL FILL_0__13458_ (
);

OR2X2 _13743_ (
    .A(_3216_),
    .B(_3215_),
    .Y(_3217_)
);

FILL FILL_0__13038_ (
);

XOR2X1 _13323_ (
    .A(_2186_),
    .B(_2863_),
    .Y(_2864_)
);

FILL FILL172520x266760 (
);

FILL FILL_1__9067_ (
);

OR2X2 _14948_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [21]),
    .Y(_3978_)
);

FILL FILL126920x0 (
);

OR2X2 _14528_ (
    .A(IRWrite_bF$buf3),
    .B(\datapath_1.PCJump [12]),
    .Y(_3758_)
);

AND2X2 _14108_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3512_)
);

FILL FILL73720x350740 (
);

FILL FILL_0__15604_ (
);

FILL FILL491720x237120 (
);

OR2X2 _18781_ (
    .A(_7684_),
    .B(_7683_),
    .Y(_7685_)
);

FILL FILL_0__18076_ (
);

OR2X2 _18361_ (
    .A(_7270_),
    .B(_7271_),
    .Y(_7272_)
);

FILL FILL390640x256880 (
);

FILL FILL_0__8597_ (
);

FILL FILL464360x172900 (
);

AND2X2 _10868_ (
    .A(_1250_),
    .B(_1249_),
    .Y(_1191_[29])
);

AND2X2 _10448_ (
    .A(_1030_),
    .B(_1029_),
    .Y(_993_[18])
);

AND2X2 _10028_ (
    .A(_810_),
    .B(_809_),
    .Y(_795_[7])
);

FILL FILL110960x54340 (
);

FILL FILL_1__12531_ (
);

FILL FILL_0__16809_ (
);

FILL FILL_0__11944_ (
);

FILL FILL_0__11104_ (
);

AND2X2 _19146_ (
    .A(_6287__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_8045_)
);

FILL FILL118560x14820 (
);

AND2X2 _14281_ (
    .A(_3633_),
    .B(_3632_),
    .Y(_3606_[13])
);

FILL FILL108680x237120 (
);

FILL FILL_1__13736_ (
);

FILL FILL_0__12729_ (
);

AND2X2 _15486_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_4440_)
);

INVX1 _15066_ (
    .A(\datapath_1.a3 [1]),
    .Y(_4054_)
);

FILL FILL_1__8758_ (
);

FILL FILL_0__16982_ (
);

FILL FILL371640x202540 (
);

FILL FILL329840x14820 (
);

FILL FILL_1__18774_ (
);

FILL FILL_0__17767_ (
);

OR2X2 _17632_ (
    .A(_6552_),
    .B(_6553_),
    .Y(_6554_)
);

FILL FILL_0__17347_ (
);

AND2X2 _17212_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_6139_)
);

FILL FILL282720x365560 (
);

FILL FILL_0__12482_ (
);

FILL FILL279680x316160 (
);

DFFSR _9974_ (
    .CLK(clk_bF$buf17),
    .D(_729_[2]),
    .Q(\datapath_1.regfile_1.regOut[12] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _9554_ (
    .A(_574_),
    .B(_573_),
    .Y(_531_[21])
);

AND2X2 _9134_ (
    .A(_354_),
    .B(_353_),
    .Y(_333_[10])
);

OR2X2 _18837_ (
    .A(_7725_),
    .B(_7740_),
    .Y(_7741_)
);

FILL FILL_0_BUFX2_insert541 (
);

AND2X2 _18417_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_7327_)
);

FILL FILL_0_BUFX2_insert543 (
);

OR2X2 _13972_ (
    .A(_3395_),
    .B(_3394_),
    .Y(_3396_)
);

FILL FILL_0__13687_ (
);

FILL FILL_0_BUFX2_insert545 (
);

OR2X2 _13552_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [21]),
    .Y(_3056_)
);

INVX1 _13132_ (
    .A(_2684_),
    .Y(\datapath_1.ALUResult [19])
);

FILL FILL_0_BUFX2_insert547 (
);

FILL FILL_0_BUFX2_insert548 (
);

FILL FILL_0_BUFX2_insert549 (
);

FILL FILL430160x44460 (
);

FILL FILL_1__15479_ (
);

FILL FILL310080x128440 (
);

OR2X2 _14757_ (
    .A(\datapath_1.rd2 [0]),
    .B(_3935__bF$buf1),
    .Y(_3871_)
);

DFFSR _14337_ (
    .CLK(clk_bF$buf62),
    .D(_3606_[1]),
    .Q(ALUOut[1]),
    .R(rst_bF$buf18),
    .S(vdd)
);

FILL FILL_0__15833_ (
);

FILL FILL_0__15413_ (
);

FILL FILL97280x34580 (
);

OR2X2 _18590_ (
    .A(_7495_),
    .B(_7496_),
    .Y(_7497_)
);

OR2X2 _18170_ (
    .A(_7076_),
    .B(_7083_),
    .Y(_7084_)
);

FILL FILL344280x281580 (
);

FILL FILL193800x316160 (
);

FILL FILL350360x222300 (
);

FILL FILL_1__17625_ (
);

OR2X2 _10677_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_1143_)
);

DFFSR _10257_ (
    .CLK(clk_bF$buf59),
    .D(_861_[27]),
    .Q(\datapath_1.regfile_1.regOut[14] [27]),
    .R(rst_bF$buf25),
    .S(vdd)
);

FILL FILL_1__12340_ (
);

OR2X2 _16903_ (
    .A(_5833_),
    .B(_5834_),
    .Y(_5835_)
);

FILL FILL_0__11333_ (
);

OR2X2 _19375_ (
    .A(_8269_),
    .B(_8262_),
    .Y(_8270_)
);

AND2X2 _14090_ (
    .A(_3352__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3497_)
);

DFFSR _8825_ (
    .CLK(clk_bF$buf1),
    .D(_135_[14]),
    .Q(\datapath_1.regfile_1.regOut[3] [14]),
    .R(rst_bF$buf38),
    .S(vdd)
);

BUFX2 _8405_ (
    .A(_1_[13]),
    .Y(memoryAddress[13])
);

FILL FILL_1__13965_ (
);

FILL FILL_0__12958_ (
);

AND2X2 _12823_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2388_)
);

FILL FILL_0__12538_ (
);

OR2X2 _12403_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .B(_2048__bF$buf0),
    .Y(_2034_)
);

AND2X2 _15295_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_4252_)
);

FILL FILL80560x330980 (
);

FILL FILL206720x207480 (
);

FILL FILL18240x88920 (
);

FILL FILL_0__16371_ (
);

FILL FILL98040x227240 (
);

AND2X2 _13608_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [2]),
    .Y(_3101_)
);

FILL FILL101080x256880 (
);

FILL FILL149720x158080 (
);

FILL FILL_0__17996_ (
);

FILL FILL255360x232180 (
);

FILL FILL_0__17576_ (
);

OR2X2 _17861_ (
    .A(_6779_),
    .B(_6772_),
    .Y(_6780_)
);

AND2X2 _17441_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_6366_)
);

OR2X2 _17021_ (
    .A(_5950_),
    .B(_5949_),
    .Y(_5951_)
);

OR2X2 _9783_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_687_)
);

FILL FILL272840x242060 (
);

OR2X2 _9363_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_467_)
);

FILL FILL_0__10604_ (
);

AND2X2 _18646_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_7552_)
);

OR2X2 _18226_ (
    .A(_7138_),
    .B(_7137_),
    .Y(_7139_)
);

FILL FILL_0__13496_ (
);

AND2X2 _13781_ (
    .A(_3084__bF$buf3),
    .B(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_3249_)
);

FILL FILL_0__13076_ (
);

OR2X2 _13361_ (
    .A(_2190_),
    .B(_2400_),
    .Y(_2900_)
);

FILL FILL79040x79040 (
);

FILL FILL76000x281580 (
);

FILL FILL23560x271700 (
);

FILL FILL53960x182780 (
);

DFFSR _14986_ (
    .CLK(clk_bF$buf20),
    .D(_3936_[5]),
    .Q(\datapath_1.mux_iord.din0 [5]),
    .R(rst_bF$buf29),
    .S(vdd)
);

AND2X2 _14566_ (
    .A(_3783_),
    .B(_3782_),
    .Y(_3738_[22])
);

OR2X2 _14146_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[1]),
    .Y(_3542_)
);

FILL FILL272080x9880 (
);

FILL FILL288800x14820 (
);

FILL FILL_0__15222_ (
);

FILL FILL257640x187720 (
);

FILL FILL255360x4940 (
);

OR2X2 _10486_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_1058__bF$buf0),
    .Y(_1056_)
);

OR2X2 _10066_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .B(_860__bF$buf1),
    .Y(_836_)
);

FILL FILL_1__17014_ (
);

FILL FILL_0__16847_ (
);

FILL FILL_0__16427_ (
);

OR2X2 _16712_ (
    .A(_5643_),
    .B(_5646_),
    .Y(_5647_)
);

FILL FILL208240x311220 (
);

FILL FILL_0__11562_ (
);

FILL FILL293360x266760 (
);

OR2X2 _19184_ (
    .A(_8080_),
    .B(_8081_),
    .Y(_8082_)
);

FILL FILL63080x271700 (
);

FILL FILL294880x4940 (
);

OR2X2 _8634_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_101_)
);

FILL FILL274360x4940 (
);

FILL FILL_1__13354_ (
);

OR2X2 _17917_ (
    .A(_6834_),
    .B(_6833_),
    .Y(_6835_)
);

INVX1 _12632_ (
    .A(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2197_)
);

FILL FILL_0__12347_ (
);

AND2X2 _12212_ (
    .A(_1926_),
    .B(_1925_),
    .Y(_1917_[4])
);

AND2X2 _9839_ (
    .A(_724_),
    .B(_723_),
    .Y(_663_[30])
);

AND2X2 _9419_ (
    .A(_504_),
    .B(_503_),
    .Y(_465_[19])
);

FILL FILL410400x187720 (
);

FILL FILL_0__16180_ (
);

FILL FILL293360x4940 (
);

FILL FILL_1__14559_ (
);

OR2X2 _13837_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [7]),
    .Y(_3291_)
);

AND2X2 _13417_ (
    .A(_2950_),
    .B(_2951_),
    .Y(_2952_)
);

FILL FILL_1__15920_ (
);

FILL FILL190000x256880 (
);

AND2X2 _17670_ (
    .A(_6591_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.rd1 [4])
);

FILL FILL_0__17385_ (
);

AND2X2 _17250_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_6177_)
);

FILL FILL228760x59280 (
);

FILL FILL255360x370500 (
);

DFFSR _9592_ (
    .CLK(clk_bF$buf39),
    .D(_531_[7]),
    .Q(\datapath_1.regfile_1.regOut[9] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

OR2X2 _9172_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .B(_398__bF$buf0),
    .Y(_380_)
);

FILL FILL19760x29640 (
);

FILL FILL_0__10833_ (
);

FILL FILL_0__10413_ (
);

AND2X2 _18875_ (
    .A(_6297__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_7778_)
);

FILL FILL_0_BUFX2_insert921 (
);

AND2X2 _18455_ (
    .A(_6211__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_7364_)
);

OR2X2 _18035_ (
    .A(_6949_),
    .B(_6950_),
    .Y(_6951_)
);

FILL FILL_0_BUFX2_insert923 (
);

AND2X2 _13590_ (
    .A(_3084__bF$buf0),
    .B(gnd),
    .Y(_3085_)
);

FILL FILL_0_BUFX2_insert925 (
);

INVX1 _13170_ (
    .A(_2697_),
    .Y(_2720_)
);

FILL FILL_0_BUFX2_insert927 (
);

FILL FILL_0_BUFX2_insert928 (
);

FILL FILL_0_BUFX2_insert929 (
);

FILL FILL_0__19111_ (
);

FILL FILL8360x138320 (
);

FILL FILL129200x182780 (
);

FILL FILL_0__11618_ (
);

AND2X2 _11903_ (
    .A(_1780_),
    .B(_1779_),
    .Y(_1719_[30])
);

OR2X2 _14795_ (
    .A(vdd),
    .B(_2_[13]),
    .Y(_3896_)
);

OR2X2 _14375_ (
    .A(vdd),
    .B(\datapath_1.Data [2]),
    .Y(_3676_)
);

FILL FILL_0__15871_ (
);

FILL FILL_0__15451_ (
);

FILL FILL143640x237120 (
);

FILL FILL_1__17243_ (
);

AND2X2 _10295_ (
    .A(_948_),
    .B(_947_),
    .Y(_927_[10])
);

AND2X2 _16941_ (
    .A(_4223__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_5873_)
);

OR2X2 _16521_ (
    .A(_5458_),
    .B(_5451_),
    .Y(_5459_)
);

FILL FILL_0__16236_ (
);

AND2X2 _16101_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_5046_)
);

FILL FILL237120x9880 (
);

FILL FILL479560x98800 (
);

OR2X2 _8863_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .B(_266__bF$buf3),
    .Y(_214_)
);

BUFX2 _8443_ (
    .A(_2_[19]),
    .Y(memoryWriteData[19])
);

FILL FILL_1__18448_ (
);

FILL FILL503880x261820 (
);

OR2X2 _17726_ (
    .A(_6645_),
    .B(_6646_),
    .Y(_6647_)
);

AND2X2 _17306_ (
    .A(_6231_),
    .B(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_6232_)
);

NAND2X1 _12861_ (
    .A(_2229_),
    .B(_2425_),
    .Y(_2426_)
);

FILL FILL_0__12576_ (
);

DFFSR _12441_ (
    .CLK(clk_bF$buf3),
    .D(_1983_[18]),
    .Q(\datapath_1.regfile_1.regOut[31] [18]),
    .R(rst_bF$buf58),
    .S(vdd)
);

FILL FILL_0__12156_ (
);

OR2X2 _12021_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_1839_)
);

FILL FILL256120x9880 (
);

FILL FILL61560x237120 (
);

OR2X2 _9648_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_617_)
);

FILL FILL177840x256880 (
);

DFFSR _9228_ (
    .CLK(clk_bF$buf108),
    .D(_333_[30]),
    .Q(\datapath_1.regfile_1.regOut[6] [30]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL384560x0 (
);

FILL FILL_0__8903_ (
);

FILL FILL118560x242060 (
);

FILL FILL_1__14368_ (
);

OR2X2 _13646_ (
    .A(_3133_),
    .B(_3130_),
    .Y(\datapath_1.mux_pcsrc.dout [7])
);

OR2X2 _13226_ (
    .A(_2420_),
    .B(_2730_),
    .Y(_2773_)
);

FILL FILL351880x172900 (
);

FILL FILL239400x4940 (
);

FILL FILL_0__14722_ (
);

FILL FILL_0__14302_ (
);

FILL FILL_0__17194_ (
);

FILL FILL_0_CLKBUF1_insert150 (
);

FILL FILL258400x4940 (
);

FILL FILL_0_CLKBUF1_insert152 (
);

FILL FILL_0__15927_ (
);

FILL FILL_0_CLKBUF1_insert154 (
);

FILL FILL_0_CLKBUF1_insert156 (
);

FILL FILL_0_CLKBUF1_insert157 (
);

FILL FILL_0__10222_ (
);

FILL FILL_0_CLKBUF1_insert158 (
);

FILL FILL_0_CLKBUF1_insert159 (
);

AND2X2 _18684_ (
    .A(_6302__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_7590_)
);

FILL FILL_0__18399_ (
);

AND2X2 _18264_ (
    .A(_6244__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_7176_)
);

FILL FILL418000x148200 (
);

FILL FILL_0__19340_ (
);

FILL FILL_1__12854_ (
);

FILL FILL_0__11847_ (
);

FILL FILL_0__9021_ (
);

OR2X2 _11712_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_1673_)
);

OR2X2 _19469_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_8348_)
);

OR2X2 _19049_ (
    .A(_7947_),
    .B(_7948_),
    .Y(_7949_)
);

FILL FILL285000x222300 (
);

AND2X2 _14184_ (
    .A(_3567_),
    .B(_3566_),
    .Y(\datapath_1.mux_wd3.dout [13])
);

OR2X2 _8919_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_251_)
);

FILL FILL431680x128440 (
);

FILL FILL175560x118560 (
);

FILL FILL262960x123500 (
);

FILL FILL_1__13219_ (
);

FILL FILL412680x286520 (
);

FILL FILL_1_BUFX2_insert470 (
);

OAI21X1 _12917_ (
    .A(_2319_),
    .B(_2324_),
    .C(_2322_),
    .Y(_2482_)
);

FILL FILL_1_BUFX2_insert472 (
);

FILL FILL329840x296400 (
);

AND2X2 _15389_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_4345_)
);

FILL FILL_1__17892_ (
);

FILL FILL348080x365560 (
);

FILL FILL120840x14820 (
);

FILL FILL_0__16885_ (
);

OR2X2 _16750_ (
    .A(_5684_),
    .B(_5683_),
    .Y(_5685_)
);

FILL FILL_0__16465_ (
);

FILL FILL_0__16045_ (
);

AND2X2 _16330_ (
    .A(_4228__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_5271_)
);

FILL FILL234840x83980 (
);

FILL FILL365560x375440 (
);

AND2X2 _8672_ (
    .A(_126_),
    .B(_125_),
    .Y(_69_[28])
);

FILL FILL254600x153140 (
);

AND2X2 _17955_ (
    .A(_6264__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_6872_)
);

OR2X2 _17535_ (
    .A(_6455_),
    .B(_6458_),
    .Y(_6459_)
);

AND2X2 _17115_ (
    .A(_4241__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_6044_)
);

XOR2X1 _12670_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2235_)
);

FILL FILL_0__12385_ (
);

OR2X2 _12250_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .B(_1982__bF$buf3),
    .Y(_1952_)
);

FILL FILL219640x316160 (
);

FILL FILL_0__18611_ (
);

FILL FILL74480x276640 (
);

OR2X2 _9877_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_794__bF$buf3),
    .Y(_730_)
);

DFFSR _9457_ (
    .CLK(clk_bF$buf93),
    .D(_465_[1]),
    .Q(\datapath_1.regfile_1.regOut[8] [1]),
    .R(rst_bF$buf41),
    .S(vdd)
);

OR2X2 _9037_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_332__bF$buf1),
    .Y(_310_)
);

FILL FILL_1__14177_ (
);

AND2X2 _13875_ (
    .A(_3316_),
    .B(_3315_),
    .Y(\datapath_1.alu_1.ALUInA [19])
);

FILL FILL150480x217360 (
);

AND2X2 _13455_ (
    .A(_2987_),
    .B(_2949_),
    .Y(_2988_)
);

INVX1 _13035_ (
    .A(_2501_),
    .Y(_2593_)
);

FILL FILL323760x237120 (
);

FILL FILL_0__14951_ (
);

FILL FILL_0__14531_ (
);

FILL FILL313120x197600 (
);

FILL FILL222680x256880 (
);

FILL FILL_0__9917_ (
);

FILL FILL_1__16743_ (
);

FILL FILL190760x311220 (
);

FILL FILL_0__15316_ (
);

AND2X2 _15601_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_4554_)
);

FILL FILL_0__10871_ (
);

FILL FILL171760x148200 (
);

FILL FILL_0__10031_ (
);

AND2X2 _18493_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_7402_)
);

FILL FILL22800x64220 (
);

AND2X2 _18073_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_6988_)
);

FILL FILL63080x44460 (
);

FILL FILL427880x251940 (
);

FILL FILL423320x54340 (
);

FILL FILL129960x74100 (
);

FILL FILL_1__17108_ (
);

FILL FILL_1__12243_ (
);

OR2X2 _16806_ (
    .A(_5739_),
    .B(_5738_),
    .Y(_5740_)
);

FILL FILL_0__9670_ (
);

OR2X2 _11941_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(_1850__bF$buf1),
    .Y(_1786_)
);

FILL FILL_0__11236_ (
);

DFFSR _11521_ (
    .CLK(clk_bF$buf16),
    .D(_1521_[1]),
    .Q(\datapath_1.regfile_1.regOut[24] [1]),
    .R(rst_bF$buf20),
    .S(vdd)
);

OR2X2 _11101_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .B(_1388__bF$buf4),
    .Y(_1366_)
);

AND2X2 _19278_ (
    .A(_6272__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_8175_)
);

OR2X2 _8728_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .B(_200__bF$buf2),
    .Y(_144_)
);

NAND2X1 _12726_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(_2290_),
    .Y(_2291_)
);

DFFSR _12306_ (
    .CLK(clk_bF$buf60),
    .D(_1917_[12]),
    .Q(\datapath_1.regfile_1.regOut[30] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

FILL FILL43320x14820 (
);

OR2X2 _15198_ (
    .A(_4155_),
    .B(_4152_),
    .Y(_4156_)
);

FILL FILL_0__13802_ (
);

FILL FILL338200x217360 (
);

FILL FILL114760x365560 (
);

FILL FILL_0__16694_ (
);

FILL FILL_0__16274_ (
);

FILL FILL256120x123500 (
);

OR2X2 _8481_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_19_)
);

FILL FILL_1__18066_ (
);

FILL FILL442320x138320 (
);

FILL FILL_0__17899_ (
);

OR2X2 _17764_ (
    .A(_6683_),
    .B(_6676_),
    .Y(_6684_)
);

FILL FILL_0__17059_ (
);

AND2X2 _17344_ (
    .A(_6219_),
    .B(_6226_),
    .Y(_6270_)
);

FILL FILL50160x192660 (
);

FILL FILL20520x88920 (
);

FILL FILL277400x330980 (
);

FILL FILL319960x360620 (
);

FILL FILL_0__18000_ (
);

AND2X2 _9686_ (
    .A(_642_),
    .B(_641_),
    .Y(_597_[22])
);

AND2X2 _9266_ (
    .A(_422_),
    .B(_421_),
    .Y(_399_[11])
);

FILL FILL_1__11514_ (
);

FILL FILL48640x74100 (
);

FILL FILL_1_CLKBUF1_insert186 (
);

FILL FILL_1_CLKBUF1_insert188 (
);

FILL FILL_0__10927_ (
);

OR2X2 _18969_ (
    .A(_7836_),
    .B(_7870_),
    .Y(_7871_)
);

OR2X2 _18549_ (
    .A(_7455_),
    .B(_7456_),
    .Y(_7457_)
);

AND2X2 _18129_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_7043_)
);

FILL FILL_0__13399_ (
);

OR2X2 _13684_ (
    .A(_3164_),
    .B(_3165_),
    .Y(_3166_)
);

XOR2X1 _13264_ (
    .A(_2222_),
    .B(_2792_),
    .Y(_2808_)
);

FILL FILL341240x93860 (
);

FILL FILL_0__19205_ (
);

FILL FILL_0__14760_ (
);

FILL FILL212800x108680 (
);

FILL FILL_1__12719_ (
);

FILL FILL_0__9306_ (
);

OR2X2 _14889_ (
    .A(\datapath_1.mux_pcsrc.dout [1]),
    .B(_4001__bF$buf0),
    .Y(_3939_)
);

DFFSR _14469_ (
    .CLK(clk_bF$buf2),
    .D(_3672_[4]),
    .Q(\datapath_1.Data [4]),
    .R(rst_bF$buf26),
    .S(vdd)
);

OR2X2 _14049_ (
    .A(_3461_),
    .B(_3460_),
    .Y(_3462_)
);

FILL FILL_0__15965_ (
);

FILL FILL_0__15545_ (
);

OR2X2 _15830_ (
    .A(_4778_),
    .B(_4777_),
    .Y(_4779_)
);

OR2X2 _15410_ (
    .A(_4365_),
    .B(_4364_),
    .Y(_4366_)
);

FILL FILL184680x187720 (
);

FILL FILL_0__10680_ (
);

FILL FILL81320x79040 (
);

FILL FILL170240x83980 (
);

FILL FILL178600x143260 (
);

DFFSR _10389_ (
    .CLK(clk_bF$buf30),
    .D(_927_[30]),
    .Q(\datapath_1.regfile_1.regOut[15] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL334400x247000 (
);

OR2X2 _16615_ (
    .A(_5551_),
    .B(_5548_),
    .Y(_5552_)
);

FILL FILL13680x311220 (
);

FILL FILL_0__11885_ (
);

AND2X2 _11750_ (
    .A(_1698_),
    .B(_1697_),
    .Y(_1653_[22])
);

FILL FILL_0__11465_ (
);

AND2X2 _11330_ (
    .A(_1478_),
    .B(_1477_),
    .Y(_1455_[11])
);

FILL FILL_0__11045_ (
);

OR2X2 _19087_ (
    .A(_7986_),
    .B(_7985_),
    .Y(_7987_)
);

DFFSR _8957_ (
    .CLK(clk_bF$buf35),
    .D(_201_[17]),
    .Q(\datapath_1.regfile_1.regOut[4] [17]),
    .R(rst_bF$buf6),
    .S(vdd)
);

AND2X2 _8537_ (
    .A(_56_),
    .B(_55_),
    .Y(_3_[26])
);

FILL FILL396720x133380 (
);

FILL FILL_1_BUFX2_insert850 (
);

NAND2X1 _12955_ (
    .A(_2354_),
    .B(_2383_),
    .Y(_2518_)
);

FILL FILL_1_BUFX2_insert852 (
);

AND2X2 _12535_ (
    .A(_2096_),
    .B(_2099_),
    .Y(_2125_)
);

OR2X2 _12115_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_1916__bF$buf2),
    .Y(_1882_)
);

FILL FILL_0__13611_ (
);

FILL FILL438520x261820 (
);

FILL FILL133760x345800 (
);

FILL FILL3800x365560 (
);

FILL FILL279680x202540 (
);

BUFX2 BUFX2_insert520 (
    .A(_3084_),
    .Y(_3084__bF$buf0)
);

BUFX2 BUFX2_insert521 (
    .A(_728_),
    .Y(_728__bF$buf4)
);

FILL FILL272840x74100 (
);

BUFX2 BUFX2_insert522 (
    .A(_728_),
    .Y(_728__bF$buf3)
);

BUFX2 BUFX2_insert523 (
    .A(_728_),
    .Y(_728__bF$buf2)
);

OR2X2 _17993_ (
    .A(_6877_),
    .B(_6909_),
    .Y(_6910_)
);

BUFX2 BUFX2_insert524 (
    .A(_728_),
    .Y(_728__bF$buf1)
);

OR2X2 _17573_ (
    .A(_6495_),
    .B(_6494_),
    .Y(_6496_)
);

BUFX2 BUFX2_insert525 (
    .A(_728_),
    .Y(_728__bF$buf0)
);

FILL FILL_0__17288_ (
);

BUFX2 BUFX2_insert526 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf113)
);

OR2X2 _17153_ (
    .A(_6080_),
    .B(_6077_),
    .Y(_6081_)
);

FILL FILL214320x212420 (
);

BUFX2 BUFX2_insert527 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf112)
);

BUFX2 BUFX2_insert528 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf111)
);

BUFX2 BUFX2_insert529 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf110)
);

FILL FILL_1__16608_ (
);

OR2X2 _9495_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_535_)
);

FILL FILL144400x217360 (
);

DFFSR _9075_ (
    .CLK(clk_bF$buf108),
    .D(_267_[6]),
    .Q(\datapath_1.regfile_1.regOut[5] [6]),
    .R(rst_bF$buf66),
    .S(vdd)
);

FILL FILL_1__11323_ (
);

FILL FILL_0__8750_ (
);

FILL FILL_0__10736_ (
);

AND2X2 _10601_ (
    .A(_1112_),
    .B(_1111_),
    .Y(_1059_[26])
);

FILL FILL_0__10316_ (
);

FILL FILL_0_BUFX2_insert41 (
);

OR2X2 _18778_ (
    .A(_7681_),
    .B(_7680_),
    .Y(_7682_)
);

FILL FILL170240x158080 (
);

FILL FILL_0_BUFX2_insert43 (
);

OR2X2 _18358_ (
    .A(_7268_),
    .B(_7265_),
    .Y(_7269_)
);

FILL FILL_0_BUFX2_insert45 (
);

FILL FILL_0_BUFX2_insert46 (
);

FILL FILL_0_BUFX2_insert47 (
);

OR2X2 _13493_ (
    .A(ALUOut[1]),
    .B(_3079__bF$buf2),
    .Y(_3017_)
);

OAI21X1 _13073_ (
    .A(_2262_),
    .B(_2376__bF$buf2),
    .C(_2628_),
    .Y(_2629_)
);

FILL FILL_0_BUFX2_insert48 (
);

FILL FILL_0_BUFX2_insert49 (
);

FILL FILL_0__19434_ (
);

FILL FILL_0__19014_ (
);

FILL FILL_1__12948_ (
);

FILL FILL_0__9955_ (
);

FILL FILL349600x212420 (
);

DFFSR _11806_ (
    .CLK(clk_bF$buf110),
    .D(_1653_[28]),
    .Q(\datapath_1.regfile_1.regOut[26] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

FILL FILL_0__9115_ (
);

AND2X2 _14698_ (
    .A(_3851_),
    .B(_3850_),
    .Y(_3804_[23])
);

AND2X2 _14278_ (
    .A(_3631_),
    .B(_3630_),
    .Y(_3606_[12])
);

FILL FILL422560x19760 (
);

FILL FILL_1__16361_ (
);

FILL FILL375440x153140 (
);

FILL FILL_0__15354_ (
);

FILL FILL280440x113620 (
);

FILL FILL447640x192660 (
);

FILL FILL_1__17566_ (
);

OR2X2 _10198_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .B(_926__bF$buf2),
    .Y(_904_)
);

FILL FILL347320x286520 (
);

FILL FILL_0__16559_ (
);

OR2X2 _16844_ (
    .A(_5775_),
    .B(_5776_),
    .Y(_5777_)
);

FILL FILL_0__16139_ (
);

OR2X2 _16424_ (
    .A(_5363_),
    .B(_5356_),
    .Y(_5364_)
);

OR2X2 _16004_ (
    .A(_4948_),
    .B(_4949_),
    .Y(_4950_)
);

FILL FILL_0__11694_ (
);

FILL FILL191520x276640 (
);

FILL FILL_0__17500_ (
);

FILL FILL364800x296400 (
);

OR2X2 _8766_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_169_)
);

OR2X2 _17629_ (
    .A(_6550_),
    .B(_6549_),
    .Y(_6551_)
);

OR2X2 _17209_ (
    .A(_6105_),
    .B(_6136_),
    .Y(_6137_)
);

FILL FILL_0__12899_ (
);

NOR2X1 _12764_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2329_)
);

AND2X2 _12344_ (
    .A(_1994_),
    .B(_1993_),
    .Y(_1983_[5])
);

FILL FILL_0__18705_ (
);

FILL FILL_0__13840_ (
);

FILL FILL_0__13420_ (
);

FILL FILL140600x247000 (
);

OR2X2 _13969_ (
    .A(_3391_),
    .B(_3392_),
    .Y(_3393_)
);

OR2X2 _13549_ (
    .A(IorD_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [20]),
    .Y(_3054_)
);

XOR2X1 _13129_ (
    .A(_2281_),
    .B(_2681_),
    .Y(_2682_)
);

FILL FILL_1__15212_ (
);

OR2X2 _14910_ (
    .A(\datapath_1.mux_pcsrc.dout [8]),
    .B(_4001__bF$buf4),
    .Y(_3953_)
);

FILL FILL_0__14205_ (
);

FILL FILL341240x227240 (
);

OR2X2 _17382_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_6308_)
);

FILL FILL345040x148200 (
);

FILL FILL_0__10965_ (
);

FILL FILL_0__10545_ (
);

OR2X2 _10830_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_1225_)
);

OR2X2 _10410_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_1005_)
);

OR2X2 _18587_ (
    .A(_7490_),
    .B(_7493_),
    .Y(_7494_)
);

AND2X2 _18167_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_7081_)
);

FILL FILL_0__9764_ (
);

AND2X2 _11615_ (
    .A(_1628_),
    .B(_1627_),
    .Y(_1587_[20])
);

FILL FILL323000x19760 (
);

AND2X2 _14087_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3494_)
);

FILL FILL388360x192660 (
);

FILL FILL117040x79040 (
);

FILL FILL_0__15583_ (
);

FILL FILL_0__15163_ (
);

FILL FILL202160x350740 (
);

FILL FILL_0__16788_ (
);

AND2X2 _16653_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_5589_)
);

FILL FILL_0__16368_ (
);

AND2X2 _16233_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_5176_)
);

FILL FILL_0__11083_ (
);

FILL FILL337440x163020 (
);

OR2X2 _8995_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .B(_332__bF$buf3),
    .Y(_282_)
);

DFFSR _8575_ (
    .CLK(clk_bF$buf91),
    .D(_3_[22]),
    .Q(\datapath_1.regfile_1.regOut[1] [22]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL328320x79040 (
);

FILL FILL_1__10403_ (
);

FILL FILL_1__13295_ (
);

AND2X2 _17858_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_6777_)
);

OR2X2 _17438_ (
    .A(_6359_),
    .B(_6362_),
    .Y(_6363_)
);

AND2X2 _17018_ (
    .A(_5948_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd2 [27])
);

NAND2X1 _12993_ (
    .A(_2476_),
    .B(_2477_),
    .Y(_2554_)
);

FILL FILL_1__19521_ (
);

FILL FILL_0__12288_ (
);

OR2X2 _12573_ (
    .A(\control_1.next [0]),
    .B(_2145_),
    .Y(_2146_)
);

OR2X2 _12153_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_1907_)
);

FILL FILL_0__18514_ (
);

FILL FILL382280x133380 (
);

FILL FILL118560x88920 (
);

FILL FILL_0__8615_ (
);

FILL FILL267520x355680 (
);

OR2X2 _13778_ (
    .A(_3246_),
    .B(_3245_),
    .Y(_3247_)
);

NOR2X1 _13358_ (
    .A(_2644_),
    .B(_2406_),
    .Y(_2897_)
);

FILL FILL_1__15861_ (
);

FILL FILL_0__14434_ (
);

FILL FILL_0__14014_ (
);

BUFX2 BUFX2_insert900 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf2 )
);

BUFX2 BUFX2_insert901 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf1 )
);

BUFX2 BUFX2_insert902 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf0 )
);

BUFX2 BUFX2_insert903 (
    .A(_4130_),
    .Y(_4130__bF$buf4)
);

BUFX2 BUFX2_insert904 (
    .A(_4130_),
    .Y(_4130__bF$buf3)
);

BUFX2 BUFX2_insert905 (
    .A(_4130_),
    .Y(_4130__bF$buf2)
);

BUFX2 BUFX2_insert906 (
    .A(_4130_),
    .Y(_4130__bF$buf1)
);

OR2X2 _17191_ (
    .A(_6118_),
    .B(_6115_),
    .Y(_6119_)
);

BUFX2 BUFX2_insert907 (
    .A(_4130_),
    .Y(_4130__bF$buf0)
);

BUFX2 BUFX2_insert908 (
    .A(_6293_),
    .Y(_6293__bF$buf4)
);

BUFX2 BUFX2_insert909 (
    .A(_6293_),
    .Y(_6293__bF$buf3)
);

FILL FILL130720x311220 (
);

FILL FILL_0__15639_ (
);

AND2X2 _15924_ (
    .A(_4177__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_4872_)
);

OR2X2 _15504_ (
    .A(_4454_),
    .B(_4457_),
    .Y(_4458_)
);

FILL FILL_0__15219_ (
);

FILL FILL_0__10354_ (
);

FILL FILL394440x360620 (
);

AND2X2 _18396_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_7306_)
);

FILL FILL211280x281580 (
);

FILL FILL_0__19472_ (
);

FILL FILL205200x64220 (
);

FILL FILL_0__19052_ (
);

FILL FILL_1__12566_ (
);

FILL FILL504640x311220 (
);

AND2X2 _16709_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_5644_)
);

FILL FILL312360x128440 (
);

FILL FILL_0__11979_ (
);

OR2X2 _11844_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_1741_)
);

FILL FILL_0__9153_ (
);

INVX2 _11424_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .Y(_1586_)
);

DFFSR _11004_ (
    .CLK(clk_bF$buf105),
    .D(_1257_[0]),
    .Q(\datapath_1.regfile_1.regOut[20] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

FILL FILL_0__12920_ (
);

FILL FILL_0__12500_ (
);

FILL FILL79800x54340 (
);

FILL FILL_0__15392_ (
);

FILL FILL346560x281580 (
);

FILL FILL265240x217360 (
);

INVX1 _12629_ (
    .A(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2194_)
);

AND2X2 _12209_ (
    .A(_1924_),
    .B(_1923_),
    .Y(_1917_[3])
);

FILL FILL_1__14712_ (
);

FILL FILL_0__13705_ (
);

FILL FILL_1__17184_ (
);

FILL FILL282720x227240 (
);

OR2X2 _16882_ (
    .A(_5813_),
    .B(_5814_),
    .Y(_5815_)
);

AND2X2 _16462_ (
    .A(_4203__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_5401_)
);

AND2X2 _16042_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .Y(_4988_)
);

FILL FILL_1__9314_ (
);

FILL FILL136040x49400 (
);

FILL FILL_1__10212_ (
);

OR2X2 _17667_ (
    .A(_6573_),
    .B(_6588_),
    .Y(_6589_)
);

OR2X2 _17247_ (
    .A(_6173_),
    .B(_6172_),
    .Y(_6174_)
);

FILL FILL410400x88920 (
);

OR2X2 _12382_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .B(_2048__bF$buf3),
    .Y(_2020_)
);

FILL FILL_0__12097_ (
);

FILL FILL_0__18743_ (
);

FILL FILL_0__18323_ (
);

DFFSR _9589_ (
    .CLK(clk_bF$buf82),
    .D(_531_[4]),
    .Q(\datapath_1.regfile_1.regOut[9] [4]),
    .R(rst_bF$buf17),
    .S(vdd)
);

OR2X2 _9169_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .B(_398__bF$buf0),
    .Y(_378_)
);

FILL FILL_0__8844_ (
);

FILL FILL_0__8424_ (
);

FILL FILL_0_BUFX2_insert890 (
);

FILL FILL_0_BUFX2_insert891 (
);

FILL FILL_0_BUFX2_insert892 (
);

FILL FILL_0_BUFX2_insert893 (
);

FILL FILL103360x256880 (
);

FILL FILL_0_BUFX2_insert894 (
);

FILL FILL_0_BUFX2_insert895 (
);

AND2X2 _13587_ (
    .A(_3081__bF$buf2),
    .B(ALUOut[0]),
    .Y(_3082_)
);

NOR2X1 _13167_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2717_)
);

FILL FILL_0_BUFX2_insert897 (
);

FILL FILL347320x49400 (
);

FILL FILL_0_BUFX2_insert899 (
);

FILL FILL_0__14663_ (
);

FILL FILL_0__14243_ (
);

FILL FILL240160x316160 (
);

FILL FILL120840x266760 (
);

FILL FILL126160x340860 (
);

FILL FILL_0__9629_ (
);

FILL FILL50920x74100 (
);

FILL FILL_1__16035_ (
);

FILL FILL_1__11170_ (
);

FILL FILL_0__15868_ (
);

OR2X2 _15733_ (
    .A(_4682_),
    .B(_4683_),
    .Y(_4684_)
);

FILL FILL_0__15028_ (
);

AND2X2 _15313_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_4270_)
);

FILL FILL481080x9880 (
);

FILL FILL_0__10163_ (
);

BUFX2 BUFX2_insert50 (
    .A(_926_),
    .Y(_926__bF$buf4)
);

BUFX2 BUFX2_insert51 (
    .A(_926_),
    .Y(_926__bF$buf3)
);

BUFX2 BUFX2_insert52 (
    .A(_926_),
    .Y(_926__bF$buf2)
);

BUFX2 BUFX2_insert53 (
    .A(_926_),
    .Y(_926__bF$buf1)
);

BUFX2 BUFX2_insert54 (
    .A(_926_),
    .Y(_926__bF$buf0)
);

BUFX2 BUFX2_insert55 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf4 )
);

BUFX2 BUFX2_insert56 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf3 )
);

BUFX2 BUFX2_insert57 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf2 )
);

BUFX2 BUFX2_insert58 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf1 )
);

BUFX2 BUFX2_insert59 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf0 )
);

FILL FILL_1__12375_ (
);

FILL FILL325280x167960 (
);

AND2X2 _16938_ (
    .A(_4146__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_5870_)
);

AND2X2 _16518_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_5456_)
);

DFFSR _11653_ (
    .CLK(clk_bF$buf83),
    .D(_1587_[4]),
    .Q(\datapath_1.regfile_1.regOut[25] [4]),
    .R(rst_bF$buf17),
    .S(vdd)
);

FILL FILL_0__11368_ (
);

OR2X2 _11233_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .B(_1454__bF$buf0),
    .Y(_1434_)
);

FILL FILL75240x326040 (
);

FILL FILL348080x251940 (
);

FILL FILL436240x98800 (
);

FILL FILL259920x187720 (
);

OR2X2 _9801_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_699_)
);

FILL FILL278160x256880 (
);

NAND2X1 _12858_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2423_)
);

DFFSR _12438_ (
    .CLK(clk_bF$buf111),
    .D(_1983_[15]),
    .Q(\datapath_1.regfile_1.regOut[31] [15]),
    .R(rst_bF$buf108),
    .S(vdd)
);

OR2X2 _12018_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_1837_)
);

FILL FILL_1__14521_ (
);

FILL FILL_1__14101_ (
);

FILL FILL_0__13934_ (
);

FILL FILL295640x266760 (
);

FILL FILL65360x271700 (
);

AND2X2 _16691_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_5627_)
);

OR2X2 _16271_ (
    .A(_5212_),
    .B(_5211_),
    .Y(_5213_)
);

FILL FILL_1__9123_ (
);

FILL FILL_1__15726_ (
);

FILL FILL265240x88920 (
);

FILL FILL_1__10021_ (
);

FILL FILL_0__14719_ (
);

AND2X2 _17896_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_6814_)
);

AND2X2 _17476_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_6400_)
);

OR2X2 _17056_ (
    .A(_5985_),
    .B(_5982_),
    .Y(_5986_)
);

DFFSR _12191_ (
    .CLK(clk_bF$buf86),
    .D(_1851_[26]),
    .Q(\datapath_1.regfile_1.regOut[29] [26]),
    .R(rst_bF$buf84),
    .S(vdd)
);

FILL FILL317680x182780 (
);

FILL FILL236360x118560 (
);

FILL FILL_0__18972_ (
);

FILL FILL_0__18552_ (
);

FILL FILL_0__18132_ (
);

AND2X2 _9398_ (
    .A(_490_),
    .B(_489_),
    .Y(_465_[12])
);

FILL FILL_1__11646_ (
);

OR2X2 _10924_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .B(_1322__bF$buf4),
    .Y(_1268_)
);

FILL FILL_0__10219_ (
);

DFFSR _10504_ (
    .CLK(clk_bF$buf97),
    .D(_993_[16]),
    .Q(\datapath_1.regfile_1.regOut[16] [16]),
    .R(rst_bF$buf84),
    .S(vdd)
);

FILL FILL110200x158080 (
);

OR2X2 _13396_ (
    .A(_2387__bF$buf0),
    .B(_2932_),
    .Y(_2933_)
);

OR2X2 _19202_ (
    .A(_8099_),
    .B(_8096_),
    .Y(_8100_)
);

FILL FILL_0__14892_ (
);

FILL FILL253080x355680 (
);

FILL FILL_0__14052_ (
);

FILL FILL458280x163020 (
);

FILL FILL67640x207480 (
);

FILL FILL_0__9438_ (
);

OR2X2 _11709_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_1671_)
);

FILL FILL_0__9018_ (
);

FILL FILL257640x370500 (
);

FILL FILL_1__16684_ (
);

AND2X2 _15962_ (
    .A(_4228__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_4909_)
);

FILL FILL_0__15677_ (
);

OR2X2 _15542_ (
    .A(_4495_),
    .B(_4492_),
    .Y(_4496_)
);

FILL FILL_0__15257_ (
);

AND2X2 _15122_ (
    .A(_4099_),
    .B(_4034_),
    .Y(_4100_)
);

FILL FILL_0__10392_ (
);

FILL FILL15200x163020 (
);

FILL FILL_0__19090_ (
);

FILL FILL498560x98800 (
);

FILL FILL_1__17049_ (
);

OR2X2 _16747_ (
    .A(_5680_),
    .B(_5681_),
    .Y(_5682_)
);

OR2X2 _16327_ (
    .A(_5267_),
    .B(_5266_),
    .Y(_5268_)
);

FILL FILL_0__11597_ (
);

AND2X2 _11882_ (
    .A(_1766_),
    .B(_1765_),
    .Y(_1719_[23])
);

FILL FILL_0__9191_ (
);

AND2X2 _11462_ (
    .A(_1546_),
    .B(_1545_),
    .Y(_1521_[12])
);

FILL FILL_0__11177_ (
);

AND2X2 _11042_ (
    .A(_1326_),
    .B(_1325_),
    .Y(_1323_[1])
);

FILL FILL_0__17823_ (
);

AND2X2 _8669_ (
    .A(_124_),
    .B(_123_),
    .Y(_69_[27])
);

DFFSR _9610_ (
    .CLK(clk_bF$buf102),
    .D(_531_[25]),
    .Q(\datapath_1.regfile_1.regOut[9] [25]),
    .R(rst_bF$buf101),
    .S(vdd)
);

FILL FILL_1__13389_ (
);

FILL FILL285000x158080 (
);

FILL FILL372400x163020 (
);

FILL FILL38000x113620 (
);

OR2X2 _12667_ (
    .A(_2229_),
    .B(_2231_),
    .Y(_2232_)
);

FILL FILL251560x311220 (
);

OR2X2 _12247_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_1982__bF$buf3),
    .Y(_1950_)
);

FILL FILL210520x9880 (
);

FILL FILL_0__13323_ (
);

OR2X2 _16080_ (
    .A(_5024_),
    .B(_5021_),
    .Y(_5025_)
);

FILL FILL249280x291460 (
);

OR2X2 _14813_ (
    .A(vdd),
    .B(_2_[19]),
    .Y(_3908_)
);

FILL FILL_0__14528_ (
);

FILL FILL_0__14108_ (
);

AND2X2 _17285_ (
    .A(_6210_),
    .B(\datapath_1.PCJump_27_bF$buf0 ),
    .Y(_6211_)
);

FILL FILL72200x360620 (
);

FILL FILL63840x237120 (
);

FILL FILL386840x311220 (
);

FILL FILL_0__18781_ (
);

FILL FILL304000x311220 (
);

FILL FILL285760x330980 (
);

FILL FILL367840x148200 (
);

FILL FILL_1__11455_ (
);

FILL FILL_0__8882_ (
);

FILL FILL_0__10868_ (
);

FILL FILL_0__10448_ (
);

AND2X2 _10733_ (
    .A(_1180_),
    .B(_1179_),
    .Y(_1125_[27])
);

FILL FILL_0__10028_ (
);

AND2X2 _10313_ (
    .A(_960_),
    .B(_959_),
    .Y(_927_[16])
);

OR2X2 _19431_ (
    .A(gnd),
    .B(_8385__bF$buf1),
    .Y(_8323_)
);

FILL FILL_0__19146_ (
);

AND2X2 _19011_ (
    .A(_6300__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_7912_)
);

FILL FILL_0__14281_ (
);

FILL FILL127680x0 (
);

DFFSR _11938_ (
    .CLK(clk_bF$buf44),
    .D(_1719_[31]),
    .Q(\datapath_1.regfile_1.regOut[27] [31]),
    .R(rst_bF$buf16),
    .S(vdd)
);

FILL FILL_0__9247_ (
);

OR2X2 _11518_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .B(_1586__bF$buf2),
    .Y(_1584_)
);

FILL FILL_1__13601_ (
);

FILL FILL503120x138320 (
);

FILL FILL370880x44460 (
);

AND2X2 _15771_ (
    .A(_4239__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_4721_)
);

FILL FILL_0__15486_ (
);

OR2X2 _15351_ (
    .A(_4300_),
    .B(_4307_),
    .Y(_4308_)
);

FILL FILL370120x212420 (
);

FILL FILL183160x59280 (
);

FILL FILL_1__17698_ (
);

OR2X2 _16976_ (
    .A(_5903_),
    .B(_5906_),
    .Y(_5907_)
);

AND2X2 _16556_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_5494_)
);

OR2X2 _16136_ (
    .A(_5076_),
    .B(_5079_),
    .Y(_5080_)
);

FILL FILL104120x143260 (
);

OR2X2 _11691_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_1659_)
);

DFFSR _11271_ (
    .CLK(clk_bF$buf24),
    .D(_1389_[9]),
    .Q(\datapath_1.regfile_1.regOut[22] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

FILL FILL230280x83980 (
);

FILL FILL_1__9408_ (
);

FILL FILL_0__17632_ (
);

FILL FILL_0__17212_ (
);

FILL FILL177840x118560 (
);

OR2X2 _8898_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_237_)
);

OR2X2 _8478_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_17_)
);

OR2X2 _12896_ (
    .A(_2460_),
    .B(_2457_),
    .Y(_2461_)
);

OR2X2 _12476_ (
    .A(\aluControl_1.inst [3]),
    .B(\aluControl_1.inst [2]),
    .Y(_2069_)
);

DFFSR _12056_ (
    .CLK(clk_bF$buf95),
    .D(_1785_[20]),
    .Q(\datapath_1.regfile_1.regOut[28] [20]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL_0__18837_ (
);

AND2X2 _18702_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_7608_)
);

FILL FILL_0__18417_ (
);

FILL FILL245480x187720 (
);

FILL FILL_0__13972_ (
);

FILL FILL_0__13552_ (
);

FILL FILL_0__13132_ (
);

FILL FILL163400x29640 (
);

FILL FILL395960x108680 (
);

FILL FILL_0__8518_ (
);

FILL FILL252320x0 (
);

FILL FILL400520x113620 (
);

DFFSR _14622_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[28]),
    .Q(\control_1.op [2]),
    .R(rst_bF$buf100),
    .S(vdd)
);

AND2X2 _14202_ (
    .A(_3579_),
    .B(_3578_),
    .Y(\datapath_1.mux_wd3.dout [19])
);

FILL FILL330600x118560 (
);

AND2X2 _17094_ (
    .A(_4146__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_6023_)
);

FILL FILL120840x88920 (
);

FILL FILL76760x276640 (
);

FILL FILL448400x242060 (
);

FILL FILL135280x207480 (
);

FILL FILL41800x64220 (
);

FILL FILL_0__18170_ (
);

FILL FILL_1__16549_ (
);

FILL FILL_1__16129_ (
);

OR2X2 _15827_ (
    .A(_4774_),
    .B(_4775_),
    .Y(_4776_)
);

OR2X2 _15407_ (
    .A(_4359_),
    .B(_4362_),
    .Y(_4363_)
);

FILL FILL503120x365560 (
);

OR2X2 _10962_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_1293_)
);

FILL FILL_0__10677_ (
);

OR2X2 _10542_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_1073_)
);

FILL FILL247000x355680 (
);

DFFSR _10122_ (
    .CLK(clk_bF$buf106),
    .D(_795_[21]),
    .Q(\datapath_1.regfile_1.regOut[13] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

OR2X2 _18299_ (
    .A(_7209_),
    .B(_7210_),
    .Y(_7211_)
);

OR2X2 _19240_ (
    .A(_8135_),
    .B(_8136_),
    .Y(_8137_)
);

FILL FILL421040x271700 (
);

FILL FILL_1__12889_ (
);

FILL FILL348840x321100 (
);

FILL FILL_0__9896_ (
);

AND2X2 _11747_ (
    .A(_1696_),
    .B(_1695_),
    .Y(_1653_[21])
);

FILL FILL_0__9056_ (
);

AND2X2 _11327_ (
    .A(_1476_),
    .B(_1475_),
    .Y(_1455_[10])
);

FILL FILL_1__13830_ (
);

FILL FILL_0__12823_ (
);

OR2X2 _15580_ (
    .A(_4531_),
    .B(_4532_),
    .Y(_4533_)
);

NAND3X1 _15160_ (
    .A(_4119_),
    .B(_4010_),
    .C(_4122_),
    .Y(_4123_)
);

FILL FILL57760x222300 (
);

FILL FILL_1__8432_ (
);

FILL FILL169480x24700 (
);

AND2X2 _16785_ (
    .A(_4181__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_5719_)
);

AND2X2 _16365_ (
    .A(_4241__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_5306_)
);

OR2X2 _11080_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .B(_1388__bF$buf4),
    .Y(_1352_)
);

FILL FILL74480x138320 (
);

FILL FILL_0__17441_ (
);

FILL FILL_0__17021_ (
);

FILL FILL_1__10955_ (
);

FILL FILL55480x296400 (
);

BUFX2 BUFX2_insert490 (
    .A(_3087_),
    .Y(_3087__bF$buf0)
);

BUFX2 BUFX2_insert491 (
    .A(_6247_),
    .Y(_6247__bF$buf4)
);

BUFX2 BUFX2_insert492 (
    .A(_6247_),
    .Y(_6247__bF$buf3)
);

BUFX2 BUFX2_insert493 (
    .A(_6247_),
    .Y(_6247__bF$buf2)
);

BUFX2 BUFX2_insert494 (
    .A(_6247_),
    .Y(_6247__bF$buf1)
);

BUFX2 BUFX2_insert495 (
    .A(_6247_),
    .Y(_6247__bF$buf0)
);

BUFX2 BUFX2_insert496 (
    .A(_4160_),
    .Y(_4160__bF$buf4)
);

BUFX2 BUFX2_insert497 (
    .A(_4160_),
    .Y(_4160__bF$buf3)
);

FILL FILL66120x14820 (
);

BUFX2 BUFX2_insert498 (
    .A(_4160_),
    .Y(_4160__bF$buf2)
);

BUFX2 BUFX2_insert499 (
    .A(_4160_),
    .Y(_4160__bF$buf1)
);

OR2X2 _12285_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_1975_)
);

FILL FILL_0__18646_ (
);

OR2X2 _18931_ (
    .A(_7832_),
    .B(_7831_),
    .Y(_7833_)
);

OR2X2 _18511_ (
    .A(_7412_),
    .B(_7419_),
    .Y(_7420_)
);

FILL FILL_0__13781_ (
);

FILL FILL_0__13361_ (
);

FILL FILL_0__8747_ (
);

FILL FILL258400x123500 (
);

FILL FILL_1__15153_ (
);

FILL FILL444600x138320 (
);

FILL FILL357960x98800 (
);

AND2X2 _14851_ (
    .A(_3933_),
    .B(_3932_),
    .Y(_3870_[31])
);

FILL FILL_0__14146_ (
);

AND2X2 _14431_ (
    .A(_3713_),
    .B(_3712_),
    .Y(_3672_[20])
);

FILL FILL76000x306280 (
);

OR2X2 _14011_ (
    .A(_3427_),
    .B(_3428_),
    .Y(_3429_)
);

FILL FILL_1__16778_ (
);

FILL FILL233320x74100 (
);

FILL FILL256120x197600 (
);

FILL FILL_1__11073_ (
);

AND2X2 _15636_ (
    .A(_4234__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_4588_)
);

OR2X2 _15216_ (
    .A(_4168_),
    .B(_4173_),
    .Y(_4174_)
);

DFFSR _10771_ (
    .CLK(clk_bF$buf16),
    .D(_1125_[25]),
    .Q(\datapath_1.regfile_1.regOut[18] [25]),
    .R(rst_bF$buf20),
    .S(vdd)
);

FILL FILL_0__10486_ (
);

FILL FILL_0__10066_ (
);

OR2X2 _10351_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .B(_992__bF$buf3),
    .Y(_986_)
);

FILL FILL_1__8908_ (
);

FILL FILL_0__16712_ (
);

FILL FILL_0__19184_ (
);

OR2X2 _11976_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_1809_)
);

OR2X2 _11556_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_1589_)
);

DFFSR _11136_ (
    .CLK(clk_bF$buf46),
    .D(_1323_[3]),
    .Q(\datapath_1.regfile_1.regOut[21] [3]),
    .R(rst_bF$buf97),
    .S(vdd)
);

FILL FILL419520x143260 (
);

FILL FILL_0__17917_ (
);

FILL FILL277400x24700 (
);

FILL FILL_0__12212_ (
);

FILL FILL263720x133380 (
);

AND2X2 _9704_ (
    .A(_654_),
    .B(_653_),
    .Y(_597_[28])
);

FILL FILL_1__14844_ (
);

FILL FILL_0__13837_ (
);

FILL FILL_0__13417_ (
);

OR2X2 _13702_ (
    .A(_3181_),
    .B(_3178_),
    .Y(\datapath_1.mux_pcsrc.dout [15])
);

FILL FILL15960x311220 (
);

AND2X2 _16594_ (
    .A(_4167__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_5531_)
);

OR2X2 _16174_ (
    .A(_5116_),
    .B(_5117_),
    .Y(_5118_)
);

FILL FILL_1__9026_ (
);

FILL FILL_0__17670_ (
);

FILL FILL_0__17250_ (
);

FILL FILL_1__10344_ (
);

OR2X2 _14907_ (
    .A(\datapath_1.mux_pcsrc.dout [7]),
    .B(_4001__bF$buf2),
    .Y(_3951_)
);

OR2X2 _17799_ (
    .A(_6685_),
    .B(_6718_),
    .Y(_6719_)
);

OR2X2 _17379_ (
    .A(_6299_),
    .B(_6304_),
    .Y(_6305_)
);

FILL FILL_1__19462_ (
);

OR2X2 _12094_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .B(_1916__bF$buf3),
    .Y(_1868_)
);

FILL FILL453720x256880 (
);

OR2X2 _18740_ (
    .A(_7631_),
    .B(_7644_),
    .Y(_7645_)
);

AND2X2 _18320_ (
    .A(_7231_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.rd1 [14])
);

FILL FILL_0__18035_ (
);

FILL FILL_0__13170_ (
);

OR2X2 _10827_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_1223_)
);

OR2X2 _10407_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_1003_)
);

FILL FILL161880x286520 (
);

NOR2X1 _13299_ (
    .A(_2423_),
    .B(_2498_),
    .Y(_2841_)
);

FILL FILL155800x242060 (
);

DFFSR _19525_ (
    .CLK(clk_bF$buf17),
    .D(_8320_[2]),
    .Q(\datapath_1.regfile_1.regOut[0] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _19105_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_8004_)
);

FILL FILL_0__14795_ (
);

OR2X2 _14660_ (
    .A(vdd),
    .B(\datapath_1.a [11]),
    .Y(_3826_)
);

INVX2 _14240_ (
    .A(vdd),
    .Y(_3671_)
);

FILL FILL36480x335920 (
);

FILL FILL_1__16167_ (
);

FILL FILL172520x158080 (
);

OR2X2 _15865_ (
    .A(_4813_),
    .B(_4782_),
    .Y(_4814_)
);

AND2X2 _15445_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_4400_)
);

NAND3X1 _15025_ (
    .A(_4013_),
    .B(\datapath_1.a3 [4]),
    .C(_4012_),
    .Y(_4014_)
);

AND2X2 _10580_ (
    .A(_1098_),
    .B(_1097_),
    .Y(_1059_[19])
);

FILL FILL_0__10295_ (
);

AND2X2 _10160_ (
    .A(_878_),
    .B(_877_),
    .Y(_861_[8])
);

FILL FILL_1__8717_ (
);

FILL FILL_0__16941_ (
);

FILL FILL_0__16521_ (
);

FILL FILL_0__16101_ (
);

FILL FILL468920x19760 (
);

DFFSR _11785_ (
    .CLK(clk_bF$buf48),
    .D(_1653_[7]),
    .Q(\datapath_1.regfile_1.regOut[26] [7]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL_1__18313_ (
);

OR2X2 _11365_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .B(_1520__bF$buf4),
    .Y(_1502_)
);

FILL FILL377720x153140 (
);

FILL FILL_0__17306_ (
);

FILL FILL282720x113620 (
);

OR2X2 _9933_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_767_)
);

OR2X2 _9513_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_547_)
);

FILL FILL117800x54340 (
);

FILL FILL293360x98800 (
);

OR2X2 _13931_ (
    .A(_3360_),
    .B(_3357_),
    .Y(\datapath_1.alu_1.ALUInB [1])
);

FILL FILL_0__13646_ (
);

FILL FILL158080x34580 (
);

FILL FILL_0__13226_ (
);

OR2X2 _13511_ (
    .A(ALUOut[7]),
    .B(_3079__bF$buf1),
    .Y(_3029_)
);

FILL FILL193800x276640 (
);

FILL FILL199120x350740 (
);

BUFX2 BUFX2_insert1050 (
    .A(_794_),
    .Y(_794__bF$buf4)
);

FILL FILL385320x365560 (
);

BUFX2 BUFX2_insert1051 (
    .A(_794_),
    .Y(_794__bF$buf3)
);

BUFX2 BUFX2_insert1052 (
    .A(_794_),
    .Y(_794__bF$buf2)
);

BUFX2 BUFX2_insert1053 (
    .A(_794_),
    .Y(_794__bF$buf1)
);

BUFX2 BUFX2_insert1054 (
    .A(_794_),
    .Y(_794__bF$buf0)
);

BUFX2 BUFX2_insert1055 (
    .A(_4203_),
    .Y(_4203__bF$buf4)
);

BUFX2 BUFX2_insert1056 (
    .A(_4203_),
    .Y(_4203__bF$buf3)
);

BUFX2 BUFX2_insert1057 (
    .A(_4203_),
    .Y(_4203__bF$buf2)
);

BUFX2 BUFX2_insert1058 (
    .A(_4203_),
    .Y(_4203__bF$buf1)
);

FILL FILL_1__15018_ (
);

BUFX2 BUFX2_insert1059 (
    .A(_4203_),
    .Y(_4203__bF$buf0)
);

FILL FILL_1__10153_ (
);

FILL FILL114000x69160 (
);

AND2X2 _14716_ (
    .A(_3863_),
    .B(_3862_),
    .Y(_3804_[29])
);

BUFX2 BUFX2_insert870 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf2 )
);

BUFX2 BUFX2_insert871 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf1 )
);

BUFX2 BUFX2_insert872 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf0 )
);

BUFX2 BUFX2_insert873 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf4 )
);

BUFX2 BUFX2_insert874 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf3 )
);

BUFX2 BUFX2_insert875 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf2 )
);

BUFX2 BUFX2_insert876 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf1 )
);

AND2X2 _17188_ (
    .A(_4234__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_6116_)
);

BUFX2 BUFX2_insert877 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf0 )
);

BUFX2 BUFX2_insert878 (
    .A(_398_),
    .Y(_398__bF$buf4)
);

BUFX2 BUFX2_insert879 (
    .A(_398_),
    .Y(_398__bF$buf3)
);

FILL FILL_0__18684_ (
);

FILL FILL_0__18264_ (
);

FILL FILL369360x34580 (
);

FILL FILL_1__11358_ (
);

FILL FILL413440x222300 (
);

FILL FILL_0__8785_ (
);

DFFSR _10636_ (
    .CLK(clk_bF$buf19),
    .D(_1059_[19]),
    .Q(\datapath_1.regfile_1.regOut[17] [19]),
    .R(rst_bF$buf19),
    .S(vdd)
);

OR2X2 _10216_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .B(_926__bF$buf3),
    .Y(_916_)
);

FILL FILL86640x0 (
);

FILL FILL116280x64220 (
);

FILL FILL_0__19469_ (
);

AND2X2 _19334_ (
    .A(_6211__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_8230_)
);

FILL FILL174040x128440 (
);

FILL FILL_0__12917_ (
);

FILL FILL152760x54340 (
);

FILL FILL_0__15389_ (
);

AND2X2 _15674_ (
    .A(_4625_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd2 [6])
);

OR2X2 _15254_ (
    .A(_4209_),
    .B(_4211_),
    .Y(_4212_)
);

FILL FILL_0__16750_ (
);

OR2X2 _16879_ (
    .A(_5808_),
    .B(_5811_),
    .Y(_5812_)
);

AND2X2 _16459_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_5398_)
);

OR2X2 _16039_ (
    .A(_4981_),
    .B(_4984_),
    .Y(_4985_)
);

FILL FILL_1__18962_ (
);

AND2X2 _11594_ (
    .A(_1614_),
    .B(_1613_),
    .Y(_1587_[13])
);

FILL FILL_1__18542_ (
);

AND2X2 _11174_ (
    .A(_1394_),
    .B(_1393_),
    .Y(_1389_[2])
);

FILL FILL318440x232180 (
);

FILL FILL_0__17535_ (
);

OR2X2 _17820_ (
    .A(_6737_),
    .B(_6738_),
    .Y(_6739_)
);

AND2X2 _17400_ (
    .A(_6296_),
    .B(_6219_),
    .Y(_6326_)
);

FILL FILL_0__17115_ (
);

FILL FILL_0__12670_ (
);

FILL FILL_0__12250_ (
);

FILL FILL152000x182780 (
);

DFFSR _9742_ (
    .CLK(clk_bF$buf110),
    .D(_597_[28]),
    .Q(\datapath_1.regfile_1.regOut[10] [28]),
    .R(rst_bF$buf74),
    .S(vdd)
);

OR2X2 _9322_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_464__bF$buf4),
    .Y(_460_)
);

INVX1 _12799_ (
    .A(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2364_)
);

OR2X2 _12379_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .B(_2048__bF$buf4),
    .Y(_2018_)
);

FILL FILL_1__19327_ (
);

FILL FILL_1__14462_ (
);

FILL FILL_1__14042_ (
);

AND2X2 _18605_ (
    .A(_6221__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_7512_)
);

FILL FILL430920x93860 (
);

FILL FILL_0__13875_ (
);

OR2X2 _13740_ (
    .A(_3212_),
    .B(_3213_),
    .Y(_3214_)
);

AND2X2 _13320_ (
    .A(_2860_),
    .B(_2200_),
    .Y(_2861_)
);

FILL FILL_1__15667_ (
);

FILL FILL_1__15247_ (
);

OR2X2 _14945_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [20]),
    .Y(_3976_)
);

OR2X2 _14525_ (
    .A(IRWrite_bF$buf3),
    .B(\datapath_1.PCJump [11]),
    .Y(_3756_)
);

OR2X2 _14105_ (
    .A(_3509_),
    .B(_3508_),
    .Y(_3510_)
);

FILL FILL_1__19080_ (
);

FILL FILL384560x133380 (
);

FILL FILL_0__18493_ (
);

FILL FILL_0__18073_ (
);

FILL FILL224200x64220 (
);

FILL FILL_0__8594_ (
);

FILL FILL462840x113620 (
);

AND2X2 _10865_ (
    .A(_1248_),
    .B(_1247_),
    .Y(_1191_[28])
);

AND2X2 _10445_ (
    .A(_1028_),
    .B(_1027_),
    .Y(_993_[17])
);

FILL FILL457520x247000 (
);

FILL FILL487920x158080 (
);

AND2X2 _10025_ (
    .A(_808_),
    .B(_807_),
    .Y(_795_[6])
);

FILL FILL418000x0 (
);

FILL FILL_0__16806_ (
);

FILL FILL_0__11941_ (
);

FILL FILL_0__19278_ (
);

OR2X2 _19143_ (
    .A(_8041_),
    .B(_8040_),
    .Y(_8042_)
);

FILL FILL373920x276640 (
);

FILL FILL_0__9379_ (
);

FILL FILL75240x54340 (
);

FILL FILL396720x360620 (
);

AND2X2 _15483_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_4437_)
);

FILL FILL_0__15198_ (
);

AND2X2 _15063_ (
    .A(_4051_),
    .B(_4047_),
    .Y(_4052_)
);

FILL FILL228000x64220 (
);

FILL FILL10640x217360 (
);

FILL FILL314640x128440 (
);

AND2X2 _16688_ (
    .A(_4236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_5624_)
);

OR2X2 _16268_ (
    .A(_5209_),
    .B(_5208_),
    .Y(_5210_)
);

FILL FILL_0__17764_ (
);

FILL FILL363280x153140 (
);

FILL FILL267520x217360 (
);

AND2X2 _9971_ (
    .A(_792_),
    .B(_791_),
    .Y(_729_[31])
);

AND2X2 _9551_ (
    .A(_572_),
    .B(_571_),
    .Y(_531_[20])
);

AND2X2 _9131_ (
    .A(_352_),
    .B(_351_),
    .Y(_333_[9])
);

FILL FILL191520x39520 (
);

DFFSR _12188_ (
    .CLK(clk_bF$buf83),
    .D(_1851_[23]),
    .Q(\datapath_1.regfile_1.regOut[29] [23]),
    .R(rst_bF$buf17),
    .S(vdd)
);

FILL FILL_1__14271_ (
);

FILL FILL380760x163020 (
);

FILL FILL_0__18549_ (
);

OR2X2 _18834_ (
    .A(_7736_),
    .B(_7737_),
    .Y(_7738_)
);

FILL FILL_0_BUFX2_insert511 (
);

FILL FILL_0__18129_ (
);

OR2X2 _18414_ (
    .A(_7323_),
    .B(_7310_),
    .Y(_7324_)
);

FILL FILL_0_BUFX2_insert512 (
);

FILL FILL_0_BUFX2_insert513 (
);

FILL FILL_0_BUFX2_insert514 (
);

FILL FILL_0_BUFX2_insert515 (
);

FILL FILL_0__13264_ (
);

FILL FILL_0_BUFX2_insert517 (
);

FILL FILL_0_BUFX2_insert519 (
);

FILL FILL196840x192660 (
);

FILL FILL_1__15896_ (
);

FILL FILL98800x306280 (
);

FILL FILL352640x296400 (
);

FILL FILL386080x103740 (
);

DFFSR _14754_ (
    .CLK(clk_bF$buf94),
    .D(_3804_[31]),
    .Q(\datapath_1.a [31]),
    .R(rst_bF$buf61),
    .S(vdd)
);

OR2X2 _14334_ (
    .A(\datapath_1.ALUResult [31]),
    .B(_3671__bF$buf4),
    .Y(_3669_)
);

FILL FILL_0__15830_ (
);

FILL FILL_0__15410_ (
);

OR2X2 _15959_ (
    .A(_4902_),
    .B(_4905_),
    .Y(_4906_)
);

AND2X2 _15539_ (
    .A(_4181__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [4]),
    .Y(_4493_)
);

AND2X2 _15119_ (
    .A(_4029_),
    .B(_4097_),
    .Y(\datapath_1.regfile_1.regEn [11])
);

OR2X2 _10674_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_1141_)
);

DFFSR _10254_ (
    .CLK(clk_bF$buf97),
    .D(_861_[24]),
    .Q(\datapath_1.regfile_1.regOut[14] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL_0__16615_ (
);

OR2X2 _16900_ (
    .A(_5830_),
    .B(_5831_),
    .Y(_5832_)
);

FILL FILL_0__11750_ (
);

FILL FILL_0__11330_ (
);

FILL FILL12160x321100 (
);

AND2X2 _19372_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_8267_)
);

FILL FILL_0__19087_ (
);

DFFSR _8822_ (
    .CLK(clk_bF$buf71),
    .D(_135_[11]),
    .Q(\datapath_1.regfile_1.regOut[3] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

BUFX2 _8402_ (
    .A(_1_[10]),
    .Y(memoryAddress[10])
);

FILL FILL_1__18827_ (
);

AND2X2 _11879_ (
    .A(_1764_),
    .B(_1763_),
    .Y(_1719_[22])
);

FILL FILL_0__9188_ (
);

FILL FILL474240x64220 (
);

AND2X2 _11459_ (
    .A(_1544_),
    .B(_1543_),
    .Y(_1521_[11])
);

FILL FILL_1__18407_ (
);

AND2X2 _11039_ (
    .A(_1324_),
    .B(_1387_),
    .Y(_1323_[0])
);

FILL FILL_0__12955_ (
);

AOI21X1 _12820_ (
    .A(_2382_),
    .B(_2384_),
    .C(_2381_),
    .Y(_2385_)
);

FILL FILL_0__12535_ (
);

OR2X2 _12400_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .B(_2048__bF$buf0),
    .Y(_2032_)
);

FILL FILL_0__12115_ (
);

FILL FILL145160x256880 (
);

AND2X2 _15292_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_4249_)
);

DFFSR _9607_ (
    .CLK(clk_bF$buf91),
    .D(_531_[22]),
    .Q(\datapath_1.regfile_1.regOut[9] [22]),
    .R(rst_bF$buf50),
    .S(vdd)
);

AND2X2 _13605_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[2]),
    .Y(_3098_)
);

AND2X2 _16497_ (
    .A(_4223__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_5436_)
);

AND2X2 _16077_ (
    .A(_4203__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_5022_)
);

FILL FILL_1__18580_ (
);

FILL FILL_1__9769_ (
);

FILL FILL39520x19760 (
);

FILL FILL_0__17153_ (
);

FILL FILL490200x360620 (
);

OR2X2 _9780_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_685_)
);

INVX2 _9360_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .Y(_530_)
);

FILL FILL380760x256880 (
);

FILL FILL63080x256880 (
);

FILL FILL386080x330980 (
);

FILL FILL468160x148200 (
);

FILL FILL297920x266760 (
);

FILL FILL_0__18778_ (
);

OR2X2 _18643_ (
    .A(_7518_),
    .B(_7549_),
    .Y(_7550_)
);

FILL FILL_0__18358_ (
);

OR2X2 _18223_ (
    .A(_7134_),
    .B(_7135_),
    .Y(_7136_)
);

FILL FILL_0__13493_ (
);

FILL FILL_0__8879_ (
);

FILL FILL_0__8459_ (
);

FILL FILL_1__12813_ (
);

FILL FILL_0__9820_ (
);

FILL FILL_0__9400_ (
);

FILL FILL_1__15285_ (
);

OR2X2 _19428_ (
    .A(gnd),
    .B(_8385__bF$buf0),
    .Y(_8321_)
);

AND2X2 _19008_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_7909_)
);

DFFSR _14983_ (
    .CLK(clk_bF$buf77),
    .D(_3936_[2]),
    .Q(\datapath_1.mux_iord.din0 [2]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL361000x217360 (
);

AND2X2 _14563_ (
    .A(_3781_),
    .B(_3780_),
    .Y(_3738_[21])
);

FILL FILL_0__14278_ (
);

INVX2 _14143_ (
    .A(MemToReg_bF$buf4),
    .Y(_3605_)
);

FILL FILL439280x232180 (
);

FILL FILL206720x79040 (
);

FILL FILL238640x118560 (
);

OR2X2 _15768_ (
    .A(_4717_),
    .B(_4710_),
    .Y(_4718_)
);

AND2X2 _15348_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_4305_)
);

FILL FILL_1__17431_ (
);

FILL FILL_0__10198_ (
);

OR2X2 _10483_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .B(_1058__bF$buf4),
    .Y(_1054_)
);

OR2X2 _10063_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .B(_860__bF$buf4),
    .Y(_834_)
);

FILL FILL_0__16004_ (
);

FILL FILL342760x360620 (
);

AND2X2 _19181_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_8079_)
);

FILL FILL69920x207480 (
);

FILL FILL434720x29640 (
);

OR2X2 _8631_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_99_)
);

OR2X2 _11688_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_1657_)
);

DFFSR _11268_ (
    .CLK(clk_bF$buf7),
    .D(_1389_[6]),
    .Q(\datapath_1.regfile_1.regOut[22] [6]),
    .R(rst_bF$buf48),
    .S(vdd)
);

FILL FILL_1__13771_ (
);

OR2X2 _17914_ (
    .A(_6830_),
    .B(_6831_),
    .Y(_6832_)
);

FILL FILL_0__17629_ (
);

FILL FILL_0__12764_ (
);

FILL FILL_0__12344_ (
);

AND2X2 _9836_ (
    .A(_722_),
    .B(_721_),
    .Y(_663_[29])
);

AND2X2 _9416_ (
    .A(_502_),
    .B(_501_),
    .Y(_465_[18])
);

FILL FILL414200x202540 (
);

FILL FILL382280x360620 (
);

FILL FILL263720x19760 (
);

FILL FILL_1__14136_ (
);

FILL FILL496280x108680 (
);

FILL FILL_0__13969_ (
);

OR2X2 _13834_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [6]),
    .Y(_3289_)
);

FILL FILL_0__13129_ (
);

INVX1 _13414_ (
    .A(_2949_),
    .Y(\datapath_1.ALUResult [2])
);

FILL FILL_0__14910_ (
);

FILL FILL_1__9158_ (
);

FILL FILL_0__17382_ (
);

FILL FILL494760x276640 (
);

FILL FILL_1__10476_ (
);

FILL FILL422560x316160 (
);

DFFSR _14619_ (
    .CLK(clk_bF$buf15),
    .D(_3738_[25]),
    .Q(\datapath_1.PCJump [27]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL253840x311220 (
);

AND2X2 _18872_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_7775_)
);

FILL FILL_0__18587_ (
);

AND2X2 _18452_ (
    .A(_6323__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_7361_)
);

OR2X2 _18032_ (
    .A(_6944_),
    .B(_6947_),
    .Y(_6948_)
);

FILL FILL340480x222300 (
);

FILL FILL_1__17907_ (
);

OR2X2 _10959_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_1291_)
);

OR2X2 _10539_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_1071_)
);

DFFSR _10119_ (
    .CLK(clk_bF$buf13),
    .D(_795_[18]),
    .Q(\datapath_1.regfile_1.regOut[13] [18]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL421800x4940 (
);

FILL FILL104120x14820 (
);

FILL FILL_0__11615_ (
);

AND2X2 _11900_ (
    .A(_1778_),
    .B(_1777_),
    .Y(_1719_[29])
);

OR2X2 _19237_ (
    .A(_8133_),
    .B(_8130_),
    .Y(_8134_)
);

OR2X2 _14792_ (
    .A(vdd),
    .B(_2_[12]),
    .Y(_3894_)
);

FILL FILL_0__14087_ (
);

OR2X2 _14372_ (
    .A(vdd),
    .B(\datapath_1.Data [1]),
    .Y(_3674_)
);

FILL FILL114000x128440 (
);

FILL FILL38760x172900 (
);

OR2X2 _15997_ (
    .A(_4941_),
    .B(_4942_),
    .Y(_4943_)
);

OR2X2 _15577_ (
    .A(_4514_),
    .B(_4529_),
    .Y(_4530_)
);

NAND2X1 _15157_ (
    .A(\datapath_1.a3 [4]),
    .B(_4013_),
    .Y(_4120_)
);

FILL FILL_1__17660_ (
);

FILL FILL500840x74100 (
);

AND2X2 _10292_ (
    .A(_946_),
    .B(_945_),
    .Y(_927_[9])
);

FILL FILL_1__8849_ (
);

FILL FILL_0__16653_ (
);

FILL FILL_0__16233_ (
);

OR2X2 _8860_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .B(_266__bF$buf3),
    .Y(_212_)
);

BUFX2 _8440_ (
    .A(_2_[16]),
    .Y(memoryWriteData[16])
);

OR2X2 _11497_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_1586__bF$buf4),
    .Y(_1570_)
);

FILL FILL505400x138320 (
);

OR2X2 _11077_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .B(_1388__bF$buf0),
    .Y(_1350_)
);

FILL FILL_1__13160_ (
);

FILL FILL_0__17858_ (
);

OR2X2 _17723_ (
    .A(_6643_),
    .B(_6640_),
    .Y(_6644_)
);

FILL FILL_0__17018_ (
);

AND2X2 _17303_ (
    .A(_6228_),
    .B(_6201_),
    .Y(_6229_)
);

FILL FILL_0__12993_ (
);

FILL FILL_0__12573_ (
);

OR2X2 _9645_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_615_)
);

DFFSR _9225_ (
    .CLK(clk_bF$buf70),
    .D(_333_[27]),
    .Q(\datapath_1.regfile_1.regOut[6] [27]),
    .R(rst_bF$buf93),
    .S(vdd)
);

FILL FILL64600x4940 (
);

FILL FILL372400x212420 (
);

FILL FILL276640x83980 (
);

FILL FILL_0__8900_ (
);

OR2X2 _18928_ (
    .A(_7829_),
    .B(_7828_),
    .Y(_7830_)
);

AND2X2 _18508_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_7417_)
);

FILL FILL_0__13778_ (
);

FILL FILL_0__13358_ (
);

AND2X2 _13643_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [7]),
    .Y(_3131_)
);

INVX1 _13223_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .Y(_2770_)
);

FILL FILL243960x266760 (
);

FILL FILL470440x192660 (
);

FILL FILL_0__17191_ (
);

FILL FILL373920x14820 (
);

FILL FILL_1__10285_ (
);

AND2X2 _14848_ (
    .A(_3931_),
    .B(_3930_),
    .Y(_3870_[30])
);

AND2X2 _14428_ (
    .A(_3711_),
    .B(_3710_),
    .Y(_3672_[19])
);

OR2X2 _14008_ (
    .A(_3426_),
    .B(_3423_),
    .Y(\datapath_1.alu_1.ALUInB [12])
);

FILL FILL370120x286520 (
);

FILL FILL_0_CLKBUF1_insert120 (
);

FILL FILL_0_CLKBUF1_insert121 (
);

FILL FILL_0_CLKBUF1_insert122 (
);

FILL FILL_0__15924_ (
);

FILL FILL_0_CLKBUF1_insert123 (
);

FILL FILL_0__15504_ (
);

FILL FILL_0_CLKBUF1_insert125 (
);

FILL FILL_0_CLKBUF1_insert127 (
);

FILL FILL_0_CLKBUF1_insert129 (
);

AND2X2 _18681_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_7587_)
);

OR2X2 _18261_ (
    .A(_7172_),
    .B(_7171_),
    .Y(_7173_)
);

FILL FILL107160x98800 (
);

FILL FILL402800x113620 (
);

DFFSR _10768_ (
    .CLK(clk_bF$buf82),
    .D(_1125_[22]),
    .Q(\datapath_1.regfile_1.regOut[18] [22]),
    .R(rst_bF$buf94),
    .S(vdd)
);

OR2X2 _10348_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .B(_992__bF$buf1),
    .Y(_984_)
);

FILL FILL370880x271700 (
);

FILL FILL_0__11424_ (
);

OR2X2 _19466_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_8346_)
);

INVX1 _19046_ (
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_7946_)
);

FILL FILL143640x88920 (
);

AND2X2 _14181_ (
    .A(_3565_),
    .B(_3564_),
    .Y(\datapath_1.mux_wd3.dout [12])
);

OR2X2 _8916_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_249_)
);

FILL FILL_1__13636_ (
);

FILL FILL465120x54340 (
);

NAND3X1 _12914_ (
    .A(_2477_),
    .B(_2476_),
    .C(_2478_),
    .Y(_2479_)
);

FILL FILL_0__12629_ (
);

FILL FILL505400x365560 (
);

FILL FILL_1_BUFX2_insert443 (
);

FILL FILL41040x64220 (
);

FILL FILL_1_BUFX2_insert445 (
);

FILL FILL_1_BUFX2_insert447 (
);

FILL FILL19000x360620 (
);

AND2X2 _15386_ (
    .A(_4230__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_4342_)
);

FILL FILL_0__16882_ (
);

FILL FILL241680x128440 (
);

FILL FILL158840x138320 (
);

FILL FILL129960x59280 (
);

FILL FILL_0__17667_ (
);

AND2X2 _17952_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_6869_)
);

FILL FILL_0__17247_ (
);

AND2X2 _17532_ (
    .A(_6323__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_6456_)
);

OR2X2 _17112_ (
    .A(_6040_),
    .B(_6033_),
    .Y(_6041_)
);

FILL FILL_0__12382_ (
);

FILL FILL186960x0 (
);

DFFSR _9874_ (
    .CLK(clk_bF$buf71),
    .D(_663_[31]),
    .Q(\datapath_1.regfile_1.regOut[11] [31]),
    .R(rst_bF$buf35),
    .S(vdd)
);

OR2X2 _9454_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .B(_530__bF$buf3),
    .Y(_528_)
);

OR2X2 _9034_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .B(_332__bF$buf4),
    .Y(_308_)
);

OR2X2 _18737_ (
    .A(_7641_),
    .B(_7640_),
    .Y(_7642_)
);

OR2X2 _18317_ (
    .A(_7213_),
    .B(_7228_),
    .Y(_7229_)
);

AND2X2 _13872_ (
    .A(_3314_),
    .B(_3313_),
    .Y(\datapath_1.alu_1.ALUInA [18])
);

FILL FILL_0__13587_ (
);

AND2X2 _13452_ (
    .A(_2714_),
    .B(_2599_),
    .Y(_2985_)
);

INVX1 _13032_ (
    .A(_2334_),
    .Y(_2590_)
);

FILL FILL62320x88920 (
);

FILL FILL389120x172900 (
);

FILL FILL_1__10094_ (
);

OR2X2 _14657_ (
    .A(vdd),
    .B(\datapath_1.a [10]),
    .Y(_3824_)
);

OR2X2 _14237_ (
    .A(\datapath_1.Data [31]),
    .B(_3605__bF$buf4),
    .Y(_3603_)
);

FILL FILL131480x4940 (
);

FILL FILL_0__15733_ (
);

FILL FILL263720x0 (
);

FILL FILL360240x163020 (
);

AND2X2 _18490_ (
    .A(_6221__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_7399_)
);

AND2X2 _18070_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_6985_)
);

FILL FILL325280x326040 (
);

FILL FILL354920x182780 (
);

FILL FILL43320x123500 (
);

FILL FILL_1__17945_ (
);

AND2X2 _10997_ (
    .A(_1316_),
    .B(_1315_),
    .Y(_1257_[29])
);

AND2X2 _10577_ (
    .A(_1096_),
    .B(_1095_),
    .Y(_1059_[18])
);

FILL FILL_1__17525_ (
);

AND2X2 _10157_ (
    .A(_876_),
    .B(_875_),
    .Y(_861_[7])
);

FILL FILL150480x4940 (
);

FILL FILL_0__16518_ (
);

OR2X2 _16803_ (
    .A(_5735_),
    .B(_5736_),
    .Y(_5737_)
);

OR2X2 _19275_ (
    .A(_8168_),
    .B(_8171_),
    .Y(_8172_)
);

FILL FILL463600x74100 (
);

OR2X2 _8725_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .B(_200__bF$buf2),
    .Y(_142_)
);

FILL FILL446120x365560 (
);

FILL FILL130720x133380 (
);

FILL FILL60040x360620 (
);

FILL FILL_1__13025_ (
);

FILL FILL287280x306280 (
);

FILL FILL463600x375440 (
);

FILL FILL_0__12858_ (
);

INVX1 _12723_ (
    .A(_2277_),
    .Y(_2288_)
);

DFFSR _12303_ (
    .CLK(clk_bF$buf113),
    .D(_1917_[9]),
    .Q(\datapath_1.regfile_1.regOut[30] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

FILL FILL_0__12018_ (
);

OR2X2 _15195_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_4153_)
);

FILL FILL108680x242060 (
);

FILL FILL_0__16271_ (
);

FILL FILL467400x296400 (
);

FILL FILL504640x133380 (
);

AND2X2 _13928_ (
    .A(_3350__bF$buf2),
    .B(_2_[1]),
    .Y(_3358_)
);

OR2X2 _13508_ (
    .A(ALUOut[6]),
    .B(_3079__bF$buf2),
    .Y(_3027_)
);

FILL FILL_0__17896_ (
);

FILL FILL_0__17476_ (
);

AND2X2 _17761_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_6681_)
);

FILL FILL_0__17056_ (
);

OR2X2 _17341_ (
    .A(_6266_),
    .B(_6261_),
    .Y(_6267_)
);

FILL FILL177080x345800 (
);

FILL FILL85880x256880 (
);

AND2X2 _9683_ (
    .A(_640_),
    .B(_639_),
    .Y(_597_[21])
);

AND2X2 _9263_ (
    .A(_420_),
    .B(_419_),
    .Y(_399_[10])
);

FILL FILL_1_CLKBUF1_insert150 (
);

FILL FILL_1_CLKBUF1_insert152 (
);

FILL FILL_1_CLKBUF1_insert154 (
);

FILL FILL317680x207480 (
);

FILL FILL_1__19268_ (
);

OR2X2 _18966_ (
    .A(_7860_),
    .B(_7867_),
    .Y(_7868_)
);

AND2X2 _18546_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_7454_)
);

AND2X2 _18126_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_7040_)
);

FILL FILL_0__13396_ (
);

OR2X2 _13681_ (
    .A(_3163_),
    .B(_3160_),
    .Y(\datapath_1.mux_pcsrc.dout [12])
);

AOI21X1 _13261_ (
    .A(_2547_),
    .B(_2805_),
    .C(_2799_),
    .Y(_2806_)
);

FILL FILL269040x281580 (
);

FILL FILL_0__11709_ (
);

OR2X2 _14886_ (
    .A(\datapath_1.mux_pcsrc.dout [0]),
    .B(_4001__bF$buf0),
    .Y(_3937_)
);

DFFSR _14466_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[1]),
    .Q(\datapath_1.Data [1]),
    .R(rst_bF$buf85),
    .S(vdd)
);

OR2X2 _14046_ (
    .A(_3457_),
    .B(_3458_),
    .Y(_3459_)
);

FILL FILL_0__15122_ (
);

DFFSR _10386_ (
    .CLK(clk_bF$buf14),
    .D(_927_[27]),
    .Q(\datapath_1.regfile_1.regOut[15] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

FILL FILL459800x177840 (
);

FILL FILL_0__16747_ (
);

AND2X2 _16612_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_5549_)
);

FILL FILL_0__16327_ (
);

FILL FILL464360x19760 (
);

FILL FILL_0__11882_ (
);

FILL FILL_0__11042_ (
);

OR2X2 _19084_ (
    .A(_7982_),
    .B(_7983_),
    .Y(_7984_)
);

FILL FILL413440x158080 (
);

FILL FILL500840x163020 (
);

DFFSR _8954_ (
    .CLK(clk_bF$buf67),
    .D(_201_[14]),
    .Q(\datapath_1.regfile_1.regOut[4] [14]),
    .R(rst_bF$buf46),
    .S(vdd)
);

AND2X2 _8534_ (
    .A(_54_),
    .B(_53_),
    .Y(_3_[25])
);

FILL FILL_1__13254_ (
);

AND2X2 _17817_ (
    .A(_6247__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_6736_)
);

FILL FILL174800x158080 (
);

OR2X2 _12952_ (
    .A(_2387__bF$buf2),
    .B(_2514_),
    .Y(_2515_)
);

FILL FILL_1_BUFX2_insert823 (
);

AND2X2 _12532_ (
    .A(_2120_),
    .B(_2121_),
    .Y(_2122_)
);

FILL FILL_0__12247_ (
);

OR2X2 _12112_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_1916__bF$buf3),
    .Y(_1880_)
);

FILL FILL_1_BUFX2_insert825 (
);

FILL FILL_1_BUFX2_insert827 (
);

FILL FILL280440x232180 (
);

FILL FILL320720x54340 (
);

DFFSR _9739_ (
    .CLK(clk_bF$buf102),
    .D(_597_[25]),
    .Q(\datapath_1.regfile_1.regOut[10] [25]),
    .R(rst_bF$buf59),
    .S(vdd)
);

OR2X2 _9319_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .B(_464__bF$buf2),
    .Y(_458_)
);

FILL FILL_0__16080_ (
);

FILL FILL180120x326040 (
);

FILL FILL190760x9880 (
);

OR2X2 _13737_ (
    .A(_3211_),
    .B(_3208_),
    .Y(\datapath_1.mux_pcsrc.dout [20])
);

AND2X2 _13317_ (
    .A(_2856_),
    .B(_2857_),
    .Y(_2858_)
);

FILL FILL468160x19760 (
);

FILL FILL_0__14813_ (
);

OR2X2 _17990_ (
    .A(_6903_),
    .B(_6906_),
    .Y(_6907_)
);

AND2X2 _17570_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_6493_)
);

AND2X2 _17150_ (
    .A(_4172__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_6078_)
);

FILL FILL434720x276640 (
);

OR2X2 _9492_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_533_)
);

DFFSR _9072_ (
    .CLK(clk_bF$buf27),
    .D(_267_[3]),
    .Q(\datapath_1.regfile_1.regOut[5] [3]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL_1__19497_ (
);

FILL FILL457520x360620 (
);

FILL FILL_0__10313_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL FILL_0_BUFX2_insert12 (
);

AND2X2 _18775_ (
    .A(_7679_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd1 [21])
);

FILL FILL_0_BUFX2_insert13 (
);

AND2X2 _18355_ (
    .A(_6289__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_7266_)
);

FILL FILL_0_BUFX2_insert15 (
);

FILL FILL_0_BUFX2_insert17 (
);

OR2X2 _13490_ (
    .A(ALUOut[0]),
    .B(_3079__bF$buf2),
    .Y(_3015_)
);

NOR2X1 _13070_ (
    .A(_2263_),
    .B(_2498_),
    .Y(_2626_)
);

FILL FILL_0_BUFX2_insert19 (
);

FILL FILL298680x301340 (
);

FILL FILL_0__19431_ (
);

FILL FILL_0__19011_ (
);

FILL FILL_1__12105_ (
);

FILL FILL_0__9952_ (
);

FILL FILL_0__9532_ (
);

FILL FILL_0__11518_ (
);

DFFSR _11803_ (
    .CLK(clk_bF$buf69),
    .D(_1653_[25]),
    .Q(\datapath_1.regfile_1.regOut[26] [25]),
    .R(rst_bF$buf79),
    .S(vdd)
);

AND2X2 _14695_ (
    .A(_3849_),
    .B(_3848_),
    .Y(_3804_[22])
);

AND2X2 _14275_ (
    .A(_3629_),
    .B(_3628_),
    .Y(_3606_[11])
);

FILL FILL122360x192660 (
);

FILL FILL_0__15771_ (
);

FILL FILL_0__15351_ (
);

FILL FILL415720x222300 (
);

OR2X2 _10195_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .B(_926__bF$buf4),
    .Y(_902_)
);

FILL FILL28120x227240 (
);

FILL FILL_0__16976_ (
);

OR2X2 _16841_ (
    .A(_5773_),
    .B(_5766_),
    .Y(_5774_)
);

FILL FILL_0__16136_ (
);

AND2X2 _16421_ (
    .A(_4217__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_5361_)
);

OR2X2 _16001_ (
    .A(_4946_),
    .B(_4943_),
    .Y(_4947_)
);

FILL FILL430920x0 (
);

OR2X2 _8763_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_167_)
);

FILL FILL176320x128440 (
);

FILL FILL3800x9880 (
);

FILL FILL40280x192660 (
);

FILL FILL_1__18348_ (
);

OR2X2 _17626_ (
    .A(_6544_),
    .B(_6547_),
    .Y(_6548_)
);

OR2X2 _17206_ (
    .A(_6130_),
    .B(_6133_),
    .Y(_6134_)
);

FILL FILL_0__12896_ (
);

FILL FILL_0__12476_ (
);

NAND2X1 _12761_ (
    .A(_2321_),
    .B(_2325_),
    .Y(_2326_)
);

FILL FILL199120x212420 (
);

AND2X2 _12341_ (
    .A(_1992_),
    .B(_1991_),
    .Y(_1983_[4])
);

AND2X2 _9968_ (
    .A(_790_),
    .B(_789_),
    .Y(_729_[30])
);

AND2X2 _9548_ (
    .A(_570_),
    .B(_569_),
    .Y(_531_[19])
);

AND2X2 _9128_ (
    .A(_350_),
    .B(_349_),
    .Y(_333_[8])
);

FILL FILL_0__8803_ (
);

FILL FILL394440x118560 (
);

FILL FILL_0_BUFX2_insert480 (
);

FILL FILL_0_BUFX2_insert482 (
);

OR2X2 _13966_ (
    .A(_3390_),
    .B(_3387_),
    .Y(\datapath_1.alu_1.ALUInB [6])
);

FILL FILL_0_BUFX2_insert484 (
);

OR2X2 _13546_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [19]),
    .Y(_3052_)
);

AND2X2 _13126_ (
    .A(_2678_),
    .B(_2460_),
    .Y(_2679_)
);

FILL FILL_0_BUFX2_insert486 (
);

FILL FILL_0_BUFX2_insert487 (
);

FILL FILL_0_BUFX2_insert488 (
);

FILL FILL_0_BUFX2_insert489 (
);

FILL FILL271320x345800 (
);

FILL FILL_0__17094_ (
);

FILL FILL155800x24700 (
);

FILL FILL_1__10188_ (
);

FILL FILL251560x133380 (
);

FILL FILL_1__16414_ (
);

FILL FILL93480x83980 (
);

FILL FILL_0__10962_ (
);

FILL FILL_0__18299_ (
);

AND2X2 _18584_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_7491_)
);

AND2X2 _18164_ (
    .A(_6326__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_7078_)
);

FILL FILL_0__19240_ (
);

FILL FILL310840x271700 (
);

FILL FILL_1__12754_ (
);

FILL FILL_0__9761_ (
);

AND2X2 _11612_ (
    .A(_1626_),
    .B(_1625_),
    .Y(_1587_[19])
);

FILL FILL_0__11327_ (
);

AND2X2 _19369_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_8264_)
);

OR2X2 _14084_ (
    .A(_3491_),
    .B(_3490_),
    .Y(_3492_)
);

FILL FILL141360x172900 (
);

FILL FILL386840x133380 (
);

DFFSR _8819_ (
    .CLK(clk_bF$buf61),
    .D(_135_[8]),
    .Q(\datapath_1.regfile_1.regOut[3] [8]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL8360x143260 (
);

FILL FILL_1__13119_ (
);

NAND2X1 _12817_ (
    .A(ALUControl[1]),
    .B(_2377_),
    .Y(_2382_)
);

FILL FILL193800x9880 (
);

FILL FILL_1__14900_ (
);

OR2X2 _15289_ (
    .A(_4194_),
    .B(_4246_),
    .Y(_4247_)
);

FILL FILL_0__16785_ (
);

AND2X2 _16650_ (
    .A(_4181__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_5586_)
);

FILL FILL_0__16365_ (
);

OR2X2 _16230_ (
    .A(_5171_),
    .B(_5172_),
    .Y(_5173_)
);

FILL FILL_0__11080_ (
);

OR2X2 _8992_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .B(_332__bF$buf2),
    .Y(_280_)
);

DFFSR _8572_ (
    .CLK(clk_bF$buf16),
    .D(_3_[19]),
    .Q(\datapath_1.regfile_1.regOut[1] [19]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL_1__18997_ (
);

AND2X2 _17855_ (
    .A(_6297__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_6774_)
);

AND2X2 _17435_ (
    .A(_6321__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_6360_)
);

OR2X2 _17015_ (
    .A(_5938_),
    .B(_5945_),
    .Y(_5946_)
);

FILL FILL230280x153140 (
);

FILL FILL112480x19760 (
);

OR2X2 _12990_ (
    .A(_2324_),
    .B(_2550_),
    .Y(_2551_)
);

OR2X2 _12570_ (
    .A(_2077_),
    .B(_2090_),
    .Y(\control_1.next [3])
);

OR2X2 _12150_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_1905_)
);

FILL FILL_0__18931_ (
);

FILL FILL_0__18511_ (
);

FILL FILL12920x217360 (
);

OR2X2 _9777_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_683_)
);

DFFSR _9357_ (
    .CLK(clk_bF$buf55),
    .D(_399_[30]),
    .Q(\datapath_1.regfile_1.regOut[7] [30]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL_1__11605_ (
);

FILL FILL_1__14077_ (
);

OR2X2 _13775_ (
    .A(_3242_),
    .B(_3243_),
    .Y(_3244_)
);

NAND3X1 _13355_ (
    .A(_2379__bF$buf1),
    .B(\datapath_1.alu_1.ALUInB [5]),
    .C(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2894_)
);

FILL FILL209000x0 (
);

FILL FILL_0__14431_ (
);

FILL FILL_0__14011_ (
);

FILL FILL411160x59280 (
);

FILL FILL_1__16643_ (
);

FILL FILL_0__15636_ (
);

AND2X2 _15921_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_4869_)
);

AND2X2 _15501_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_4455_)
);

FILL FILL_0__15216_ (
);

FILL FILL_0__10351_ (
);

AND2X2 _18393_ (
    .A(_6221__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_7303_)
);

FILL FILL37240x296400 (
);

FILL FILL424080x197600 (
);

AND2X2 _16706_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_5641_)
);

FILL FILL388360x103740 (
);

FILL FILL_0__9570_ (
);

FILL FILL_0__11556_ (
);

FILL FILL_0__9150_ (
);

OR2X2 _11841_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_1739_)
);

DFFSR _11421_ (
    .CLK(clk_bF$buf108),
    .D(_1455_[30]),
    .Q(\datapath_1.regfile_1.regOut[23] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

OR2X2 _11001_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_1319_)
);

OR2X2 _19178_ (
    .A(_8075_),
    .B(_8074_),
    .Y(_8076_)
);

OR2X2 _8628_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_97_)
);

FILL FILL88160x113620 (
);

FILL FILL262200x143260 (
);

FILL FILL291080x271700 (
);

NAND2X1 _12626_ (
    .A(_2189_),
    .B(_2190_),
    .Y(_2191_)
);

AND2X2 _12206_ (
    .A(_1922_),
    .B(_1921_),
    .Y(_1917_[2])
);

FILL FILL334400x182780 (
);

INVX1 _15098_ (
    .A(_4080_),
    .Y(_4081_)
);

FILL FILL_0__13702_ (
);

FILL FILL14440x321100 (
);

FILL FILL_0__16594_ (
);

FILL FILL_0__16174_ (
);

FILL FILL504640x247000 (
);

FILL FILL_1__18386_ (
);

OR2X2 _17664_ (
    .A(_6585_),
    .B(_6584_),
    .Y(_6586_)
);

OR2X2 _17244_ (
    .A(_6169_),
    .B(_6170_),
    .Y(_6171_)
);

FILL FILL117040x345800 (
);

DFFSR _9586_ (
    .CLK(clk_bF$buf22),
    .D(_531_[1]),
    .Q(\datapath_1.regfile_1.regOut[9] [1]),
    .R(rst_bF$buf7),
    .S(vdd)
);

OR2X2 _9166_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .B(_398__bF$buf2),
    .Y(_376_)
);

FILL FILL_0__10827_ (
);

FILL FILL_0__10407_ (
);

FILL FILL315400x44460 (
);

OR2X2 _18869_ (
    .A(_7771_),
    .B(_7758_),
    .Y(_7772_)
);

FILL FILL_0_BUFX2_insert860 (
);

OR2X2 _18449_ (
    .A(_7324_),
    .B(_7358_),
    .Y(_7359_)
);

FILL FILL_0_BUFX2_insert862 (
);

AND2X2 _18029_ (
    .A(_6287__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_6945_)
);

FILL FILL205960x64220 (
);

FILL FILL_0_BUFX2_insert864 (
);

AND2X2 _13584_ (
    .A(_3077_),
    .B(_3076_),
    .Y(_1_[31])
);

FILL FILL_0__13299_ (
);

FILL FILL_0_BUFX2_insert866 (
);

INVX1 _13164_ (
    .A(_2714_),
    .Y(\datapath_1.ALUResult [17])
);

FILL FILL_0_BUFX2_insert867 (
);

FILL FILL_0_BUFX2_insert868 (
);

FILL FILL_0_BUFX2_insert869 (
);

FILL FILL367080x123500 (
);

FILL FILL_0__19105_ (
);

FILL FILL_0__14240_ (
);

FILL FILL_1__12619_ (
);

FILL FILL202160x79040 (
);

OR2X2 _14789_ (
    .A(vdd),
    .B(_2_[11]),
    .Y(_3892_)
);

INVX2 _14369_ (
    .A(vdd),
    .Y(_3737_)
);

FILL FILL_0__15865_ (
);

FILL FILL_0__15445_ (
);

OR2X2 _15730_ (
    .A(_4680_),
    .B(_4679_),
    .Y(_4681_)
);

FILL FILL144400x34580 (
);

AND2X2 _15310_ (
    .A(_4160__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_4267_)
);

FILL FILL_0__10580_ (
);

FILL FILL_0__10160_ (
);

BUFX2 BUFX2_insert20 (
    .A(_6216_),
    .Y(_6216__bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .A(_6216_),
    .Y(_6216__bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .A(_6216_),
    .Y(_6216__bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .A(_6216_),
    .Y(_6216__bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .A(_6216_),
    .Y(_6216__bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf4 )
);

BUFX2 BUFX2_insert26 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf3 )
);

BUFX2 BUFX2_insert27 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf2 )
);

BUFX2 BUFX2_insert28 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf1 )
);

BUFX2 BUFX2_insert29 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf0 )
);

FILL FILL477280x59280 (
);

AND2X2 _10289_ (
    .A(_944_),
    .B(_943_),
    .Y(_927_[8])
);

OR2X2 _16935_ (
    .A(_5863_),
    .B(_5866_),
    .Y(_5867_)
);

AND2X2 _16515_ (
    .A(_4154__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_5453_)
);

FILL FILL505400x251940 (
);

DFFSR _11650_ (
    .CLK(clk_bF$buf67),
    .D(_1587_[1]),
    .Q(\datapath_1.regfile_1.regOut[25] [1]),
    .R(rst_bF$buf7),
    .S(vdd)
);

FILL FILL_0__11365_ (
);

OR2X2 _11230_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .B(_1454__bF$buf2),
    .Y(_1432_)
);

OR2X2 _8857_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_266__bF$buf4),
    .Y(_210_)
);

BUFX2 _8437_ (
    .A(_2_[13]),
    .Y(memoryWriteData[13])
);

FILL FILL126160x276640 (
);

FILL FILL_1__13577_ (
);

XOR2X1 _12855_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2420_)
);

DFFSR _12435_ (
    .CLK(clk_bF$buf28),
    .D(_1983_[12]),
    .Q(\datapath_1.regfile_1.regOut[31] [12]),
    .R(rst_bF$buf0),
    .S(vdd)
);

FILL FILL350360x44460 (
);

OR2X2 _12015_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_1835_)
);

FILL FILL292600x192660 (
);

FILL FILL282720x19760 (
);

FILL FILL_0__13511_ (
);

FILL FILL_1__8599_ (
);

FILL FILL475760x158080 (
);

FILL FILL_1__9960_ (
);

FILL FILL_0__14716_ (
);

OR2X2 _17893_ (
    .A(_6807_),
    .B(_6810_),
    .Y(_6811_)
);

FILL FILL449160x9880 (
);

OR2X2 _17473_ (
    .A(_6366_),
    .B(_6397_),
    .Y(_6398_)
);

FILL FILL_0__17188_ (
);

AND2X2 _17053_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_5983_)
);

FILL FILL38000x232180 (
);

FILL FILL101840x148200 (
);

FILL FILL330600x14820 (
);

FILL FILL384560x360620 (
);

AND2X2 _9395_ (
    .A(_488_),
    .B(_487_),
    .Y(_465_[11])
);

FILL FILL_1__16508_ (
);

FILL FILL498560x108680 (
);

FILL FILL_0__8650_ (
);

OR2X2 _10921_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .B(_1322__bF$buf2),
    .Y(_1266_)
);

DFFSR _10501_ (
    .CLK(clk_bF$buf47),
    .D(_993_[13]),
    .Q(\datapath_1.regfile_1.regOut[16] [13]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL_0__10216_ (
);

AND2X2 _18678_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_7584_)
);

OR2X2 _18258_ (
    .A(_7169_),
    .B(_7168_),
    .Y(_7170_)
);

FILL FILL410400x355680 (
);

FILL FILL505400x24700 (
);

NOR2X1 _13393_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2930_)
);

FILL FILL_0__19334_ (
);

FILL FILL93480x261820 (
);

FILL FILL_1__12008_ (
);

FILL FILL424840x316160 (
);

FILL FILL_0__9435_ (
);

OR2X2 _11706_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_1669_)
);

DFFSR _14598_ (
    .CLK(clk_bF$buf2),
    .D(_3738_[4]),
    .Q(\aluControl_1.inst [4]),
    .R(rst_bF$buf33),
    .S(vdd)
);

AND2X2 _14178_ (
    .A(_3563_),
    .B(_3562_),
    .Y(\datapath_1.mux_wd3.dout [11])
);

FILL FILL_0__15254_ (
);

FILL FILL_1__17466_ (
);

OR2X2 _10098_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_857_)
);

OR2X2 _16744_ (
    .A(_5671_),
    .B(_5678_),
    .Y(_5679_)
);

FILL FILL_0__16459_ (
);

FILL FILL376200x256880 (
);

FILL FILL_0__16039_ (
);

OR2X2 _16324_ (
    .A(_5264_),
    .B(_5263_),
    .Y(_5265_)
);

FILL FILL_0__11174_ (
);

FILL FILL_0__17400_ (
);

AND2X2 _8666_ (
    .A(_122_),
    .B(_121_),
    .Y(_69_[26])
);

FILL FILL399000x340860 (
);

OR2X2 _17949_ (
    .A(_6864_),
    .B(_6865_),
    .Y(_6866_)
);

AND2X2 _17529_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_6453_)
);

AND2X2 _17109_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_6038_)
);

FILL FILL_0__12799_ (
);

XOR2X1 _12664_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2229_)
);

FILL FILL_0__12379_ (
);

FILL FILL480320x177840 (
);

FILL FILL339720x74100 (
);

OR2X2 _12244_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .B(_1982__bF$buf1),
    .Y(_1948_)
);

FILL FILL_0__18605_ (
);

FILL FILL_0__13740_ (
);

AND2X2 _13869_ (
    .A(_3312_),
    .B(_3311_),
    .Y(\datapath_1.alu_1.ALUInA [17])
);

AND2X2 _13449_ (
    .A(_2981_),
    .B(_2974_),
    .Y(_2982_)
);

INVX1 _13029_ (
    .A(_2587_),
    .Y(\datapath_1.ALUResult [25])
);

FILL FILL_1__15532_ (
);

FILL FILL_1__15112_ (
);

FILL FILL_0__14945_ (
);

OR2X2 _14810_ (
    .A(vdd),
    .B(_2_[18]),
    .Y(_3906_)
);

FILL FILL_0__14525_ (
);

FILL FILL_0__14105_ (
);

FILL FILL357200x202540 (
);

INVX1 _17282_ (
    .A(\datapath_1.PCJump [25]),
    .Y(_6208_)
);

FILL FILL503880x108680 (
);

FILL FILL_0__10445_ (
);

AND2X2 _10730_ (
    .A(_1178_),
    .B(_1177_),
    .Y(_1125_[26])
);

AND2X2 _10310_ (
    .A(_958_),
    .B(_957_),
    .Y(_927_[15])
);

FILL FILL_0__10025_ (
);

OR2X2 _18487_ (
    .A(_7394_),
    .B(_7395_),
    .Y(_7396_)
);

OR2X2 _18067_ (
    .A(_6980_),
    .B(_6981_),
    .Y(_6982_)
);

FILL FILL294880x0 (
);

FILL FILL_0__9664_ (
);

DFFSR _11935_ (
    .CLK(clk_bF$buf25),
    .D(_1719_[28]),
    .Q(\datapath_1.regfile_1.regOut[27] [28]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL_0__9244_ (
);

OR2X2 _11515_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .B(_1586__bF$buf1),
    .Y(_1582_)
);

FILL FILL372400x286520 (
);

FILL FILL_0__15483_ (
);

FILL FILL_0__15063_ (
);

FILL FILL386840x247000 (
);

FILL FILL69160x247000 (
);

FILL FILL26600x143260 (
);

FILL FILL_1__14803_ (
);

FILL FILL_1_BUFX2_insert80 (
);

FILL FILL_1_BUFX2_insert88 (
);

FILL FILL_0__16688_ (
);

AND2X2 _16973_ (
    .A(_4230__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_5904_)
);

AND2X2 _16553_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_5491_)
);

AND2X2 _16133_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_5077_)
);

OR2X2 _8895_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_235_)
);

OR2X2 _8475_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_15_)
);

FILL FILL421800x350740 (
);

FILL FILL_1__13195_ (
);

FILL FILL380000x83980 (
);

AND2X2 _17758_ (
    .A(_6206__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_6678_)
);

AND2X2 _17338_ (
    .A(_6231_),
    .B(_6201_),
    .Y(_6264_)
);

NOR2X1 _12893_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2458_)
);

OR2X2 _12473_ (
    .A(_2065_),
    .B(_2062_),
    .Y(_2066_)
);

DFFSR _12053_ (
    .CLK(clk_bF$buf53),
    .D(_1785_[17]),
    .Q(\datapath_1.regfile_1.regOut[28] [17]),
    .R(rst_bF$buf111),
    .S(vdd)
);

FILL FILL_0__18414_ (
);

FILL FILL243960x128440 (
);

FILL FILL_0__8935_ (
);

FILL FILL224960x286520 (
);

FILL FILL_0__8515_ (
);

AND2X2 _13678_ (
    .A(_3087__bF$buf0),
    .B(\datapath_1.ALUResult [12]),
    .Y(_3161_)
);

OR2X2 _13258_ (
    .A(_2222_),
    .B(_2802_),
    .Y(_2803_)
);

FILL FILL_1__15761_ (
);

FILL FILL_0__14334_ (
);

AND2X2 _17091_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_6020_)
);

FILL FILL387600x251940 (
);

FILL FILL123120x108680 (
);

FILL FILL210520x113620 (
);

FILL FILL9120x261820 (
);

FILL FILL_0__15959_ (
);

FILL FILL_0__15539_ (
);

OR2X2 _15824_ (
    .A(_4769_),
    .B(_4772_),
    .Y(_4773_)
);

FILL FILL_0__15119_ (
);

AND2X2 _15404_ (
    .A(_4234__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_4360_)
);

OR2X2 _18296_ (
    .A(_7206_),
    .B(_7207_),
    .Y(_7208_)
);

FILL FILL140600x118560 (
);

FILL FILL_0__16900_ (
);

FILL FILL_0__19372_ (
);

FILL FILL395960x365560 (
);

FILL FILL_1__12466_ (
);

FILL FILL78280x365560 (
);

AND2X2 _16609_ (
    .A(_4214__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_5546_)
);

FILL FILL345040x153140 (
);

FILL FILL_0__9893_ (
);

FILL FILL_0__11459_ (
);

AND2X2 _11744_ (
    .A(_1694_),
    .B(_1693_),
    .Y(_1653_[20])
);

AND2X2 _11324_ (
    .A(_1474_),
    .B(_1473_),
    .Y(_1455_[9])
);

FILL FILL275120x74100 (
);

FILL FILL104880x251940 (
);

FILL FILL_0__12820_ (
);

FILL FILL_0__12400_ (
);

FILL FILL_0__15292_ (
);

FILL FILL_1_BUFX2_insert790 (
);

OR2X2 _12949_ (
    .A(_2359_),
    .B(_2484_),
    .Y(_2512_)
);

INVX1 _12529_ (
    .A(\control_1.op [4]),
    .Y(_2119_)
);

FILL FILL45600x123500 (
);

OR2X2 _12109_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_1916__bF$buf4),
    .Y(_1878_)
);

FILL FILL_1_BUFX2_insert799 (
);

FILL FILL_0__13605_ (
);

FILL FILL_1__17084_ (
);

AND2X2 _16782_ (
    .A(_4177__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_5716_)
);

FILL FILL_0__16077_ (
);

AND2X2 _16362_ (
    .A(_4225__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_5303_)
);

FILL FILL233320x59280 (
);

FILL FILL497800x163020 (
);

FILL FILL289560x306280 (
);

BUFX2 BUFX2_insert460 (
    .A(_4225_),
    .Y(_4225__bF$buf0)
);

BUFX2 BUFX2_insert461 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf4 )
);

BUFX2 BUFX2_insert462 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf3 )
);

BUFX2 BUFX2_insert463 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf2 )
);

AND2X2 _17987_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_6904_)
);

BUFX2 BUFX2_insert464 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf1 )
);

OR2X2 _17567_ (
    .A(_6486_),
    .B(_6489_),
    .Y(_6490_)
);

BUFX2 BUFX2_insert465 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf0 )
);

BUFX2 BUFX2_insert466 (
    .A(_1388_),
    .Y(_1388__bF$buf4)
);

AND2X2 _17147_ (
    .A(_4135__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_6075_)
);

FILL FILL275880x330980 (
);

BUFX2 BUFX2_insert467 (
    .A(_1388_),
    .Y(_1388__bF$buf3)
);

BUFX2 BUFX2_insert468 (
    .A(_1388_),
    .Y(_1388__bF$buf2)
);

BUFX2 BUFX2_insert469 (
    .A(_1388_),
    .Y(_1388__bF$buf1)
);

OR2X2 _12282_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_1973_)
);

FILL FILL_0__18223_ (
);

FILL FILL224200x316160 (
);

INVX2 _9489_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .Y(_596_)
);

DFFSR _9069_ (
    .CLK(clk_bF$buf105),
    .D(_267_[0]),
    .Q(\datapath_1.regfile_1.regOut[5] [0]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL60800x19760 (
);

FILL FILL480320x98800 (
);

FILL FILL_1__11737_ (
);

AND2X2 _13487_ (
    .A(_3014_),
    .B(_3013_),
    .Y(\datapath_1.a3 [4])
);

INVX1 _13067_ (
    .A(_2623_),
    .Y(\datapath_1.ALUResult [23])
);

FILL FILL179360x345800 (
);

FILL FILL_0__14563_ (
);

FILL FILL_0__14143_ (
);

FILL FILL_0__9529_ (
);

FILL FILL237120x128440 (
);

FILL FILL_0__9109_ (
);

FILL FILL442320x306280 (
);

FILL FILL273600x301340 (
);

FILL FILL_1__11490_ (
);

FILL FILL309320x167960 (
);

FILL FILL_0__15768_ (
);

AND2X2 _15633_ (
    .A(_4203__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_4585_)
);

AND2X2 _15213_ (
    .A(_4170_),
    .B(\datapath_1.PCJump [21]),
    .Y(_4171_)
);

FILL FILL290320x217360 (
);

FILL FILL131480x83980 (
);

FILL FILL_1__12695_ (
);

AND2X2 _16838_ (
    .A(_4225__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_5771_)
);

AND2X2 _16418_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_5358_)
);

OR2X2 _11973_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_1807_)
);

FILL FILL_0__11688_ (
);

FILL FILL_1__18921_ (
);

FILL FILL_0__9282_ (
);

INVX2 _11553_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .Y(_1652_)
);

DFFSR _11133_ (
    .CLK(clk_bF$buf99),
    .D(_1323_[0]),
    .Q(\datapath_1.regfile_1.regOut[21] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL268280x326040 (
);

FILL FILL_0__17914_ (
);

FILL FILL66880x14820 (
);

AND2X2 _9701_ (
    .A(_652_),
    .B(_651_),
    .Y(_597_[27])
);

INVX1 _12758_ (
    .A(_2322_),
    .Y(_2323_)
);

AND2X2 _12338_ (
    .A(_1990_),
    .B(_1989_),
    .Y(_1983_[3])
);

FILL FILL_1__14001_ (
);

FILL FILL_0__13834_ (
);

FILL FILL12160x143260 (
);

OR2X2 _16591_ (
    .A(_5526_),
    .B(_5527_),
    .Y(_5528_)
);

OR2X2 _16171_ (
    .A(_5114_),
    .B(_5113_),
    .Y(_5115_)
);

FILL FILL239400x39520 (
);

FILL FILL_1__15626_ (
);

FILL FILL389880x350740 (
);

OR2X2 _14904_ (
    .A(\datapath_1.mux_pcsrc.dout [6]),
    .B(_4001__bF$buf2),
    .Y(_3949_)
);

FILL FILL282720x232180 (
);

OR2X2 _17796_ (
    .A(_6715_),
    .B(_6708_),
    .Y(_6716_)
);

AND2X2 _17376_ (
    .A(_6246_),
    .B(\datapath_1.PCJump_27_bF$buf1 ),
    .Y(_6302_)
);

OR2X2 _12091_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .B(_1916__bF$buf2),
    .Y(_1866_)
);

FILL FILL129960x222300 (
);

FILL FILL_0__18872_ (
);

FILL FILL_0__18452_ (
);

OR2X2 _9298_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .B(_464__bF$buf4),
    .Y(_444_)
);

FILL FILL_1__11126_ (
);

FILL FILL_0__8973_ (
);

FILL FILL_0__10959_ (
);

OR2X2 _10824_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_1221_)
);

FILL FILL_0__10539_ (
);

OR2X2 _10404_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_1001_)
);

FILL FILL52440x103740 (
);

OR2X2 _13296_ (
    .A(_2424_),
    .B(_2376__bF$buf0),
    .Y(_2838_)
);

FILL FILL_0__11900_ (
);

AND2X2 _19522_ (
    .A(_8383_),
    .B(_8382_),
    .Y(_8320_[31])
);

FILL FILL_0__19237_ (
);

AND2X2 _19102_ (
    .A(_6216__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_8001_)
);

FILL FILL_0__14372_ (
);

AND2X2 _11609_ (
    .A(_1624_),
    .B(_1623_),
    .Y(_1587_[18])
);

FILL FILL350360x167960 (
);

FILL FILL50920x271700 (
);

FILL FILL_1__16584_ (
);

OR2X2 _15862_ (
    .A(_4807_),
    .B(_4810_),
    .Y(_4811_)
);

FILL FILL_0__15577_ (
);

FILL FILL_0__15157_ (
);

AND2X2 _15442_ (
    .A(_4146__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [3]),
    .Y(_4397_)
);

OR2X2 _15022_ (
    .A(_4010_),
    .B(_4009_),
    .Y(_4011_)
);

FILL FILL218120x301340 (
);

FILL FILL107160x182780 (
);

OR2X2 _16647_ (
    .A(_5582_),
    .B(_5581_),
    .Y(_5583_)
);

OR2X2 _16227_ (
    .A(_5169_),
    .B(_5168_),
    .Y(_5170_)
);

DFFSR _11782_ (
    .CLK(clk_bF$buf24),
    .D(_1653_[4]),
    .Q(\datapath_1.regfile_1.regOut[26] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL_0__11497_ (
);

FILL FILL_0__11077_ (
);

OR2X2 _11362_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .B(_1520__bF$buf3),
    .Y(_1500_)
);

FILL FILL_0__17723_ (
);

FILL FILL26600x306280 (
);

OR2X2 _8989_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .B(_332__bF$buf3),
    .Y(_278_)
);

DFFSR _8569_ (
    .CLK(clk_bF$buf107),
    .D(_3_[16]),
    .Q(\datapath_1.regfile_1.regOut[1] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

FILL FILL_1__10817_ (
);

FILL FILL12920x330980 (
);

FILL FILL130720x74100 (
);

OR2X2 _9930_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_765_)
);

OR2X2 _9510_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_545_)
);

INVX1 _12987_ (
    .A(_2376__bF$buf3),
    .Y(_2548_)
);

OR2X2 _12567_ (
    .A(_2084_),
    .B(_2087_),
    .Y(_2088_)
);

OR2X2 _12147_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_1903_)
);

FILL FILL_1__14650_ (
);

FILL FILL_0__18928_ (
);

FILL FILL_0_BUFX2_insert101 (
);

FILL FILL_0_BUFX2_insert103 (
);

FILL FILL_0__13643_ (
);

FILL FILL_0__13223_ (
);

FILL FILL_0_BUFX2_insert105 (
);

FILL FILL_0_BUFX2_insert107 (
);

FILL FILL_0_BUFX2_insert108 (
);

FILL FILL_0_BUFX2_insert109 (
);

FILL FILL379240x242060 (
);

FILL FILL_0__8609_ (
);

FILL FILL178600x128440 (
);

BUFX2 BUFX2_insert1020 (
    .A(_530_),
    .Y(_530__bF$buf4)
);

BUFX2 BUFX2_insert1021 (
    .A(_530_),
    .Y(_530__bF$buf3)
);

BUFX2 BUFX2_insert1022 (
    .A(_530_),
    .Y(_530__bF$buf2)
);

BUFX2 BUFX2_insert1023 (
    .A(_530_),
    .Y(_530__bF$buf1)
);

FILL FILL42560x192660 (
);

BUFX2 BUFX2_insert1024 (
    .A(_530_),
    .Y(_530__bF$buf0)
);

BUFX2 BUFX2_insert1025 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf4 )
);

BUFX2 BUFX2_insert1026 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf3 )
);

FILL FILL284240x202540 (
);

BUFX2 BUFX2_insert1027 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf2 )
);

BUFX2 BUFX2_insert1028 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf1 )
);

BUFX2 BUFX2_insert1029 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf0 )
);

FILL FILL382280x54340 (
);

FILL FILL_0__14848_ (
);

AND2X2 _14713_ (
    .A(_3861_),
    .B(_3860_),
    .Y(_3804_[28])
);

FILL FILL_0__14008_ (
);

BUFX2 BUFX2_insert840 (
    .A(_134_),
    .Y(_134__bF$buf2)
);

BUFX2 BUFX2_insert841 (
    .A(_134_),
    .Y(_134__bF$buf1)
);

BUFX2 BUFX2_insert842 (
    .A(_134_),
    .Y(_134__bF$buf0)
);

BUFX2 BUFX2_insert843 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf4 )
);

BUFX2 BUFX2_insert844 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf3 )
);

BUFX2 BUFX2_insert845 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf2 )
);

BUFX2 BUFX2_insert846 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf1 )
);

AND2X2 _17185_ (
    .A(_4208__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_6113_)
);

BUFX2 BUFX2_insert847 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf0 )
);

BUFX2 BUFX2_insert848 (
    .A(_6317_),
    .Y(_6317__bF$buf4)
);

FILL FILL134520x74100 (
);

BUFX2 BUFX2_insert849 (
    .A(_6317_),
    .Y(_6317__bF$buf3)
);

FILL FILL151240x24700 (
);

FILL FILL279680x321100 (
);

OR2X2 _15918_ (
    .A(_4865_),
    .B(_4864_),
    .Y(_4866_)
);

FILL FILL_0__8782_ (
);

FILL FILL_0__10348_ (
);

DFFSR _10633_ (
    .CLK(clk_bF$buf53),
    .D(_1059_[16]),
    .Q(\datapath_1.regfile_1.regOut[17] [16]),
    .R(rst_bF$buf111),
    .S(vdd)
);

OR2X2 _10213_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .B(_926__bF$buf3),
    .Y(_914_)
);

FILL FILL364800x9880 (
);

FILL FILL_0__19466_ (
);

FILL FILL_0__19046_ (
);

AND2X2 _19331_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_8227_)
);

FILL FILL_0__14181_ (
);

FILL FILL_0__9567_ (
);

OR2X2 _11838_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_1737_)
);

FILL FILL253840x133380 (
);

DFFSR _11418_ (
    .CLK(clk_bF$buf39),
    .D(_1455_[27]),
    .Q(\datapath_1.regfile_1.regOut[23] [27]),
    .R(rst_bF$buf69),
    .S(vdd)
);

FILL FILL_1__13501_ (
);

FILL FILL155040x24700 (
);

FILL FILL208240x256880 (
);

OR2X2 _15671_ (
    .A(_4622_),
    .B(_4615_),
    .Y(_4623_)
);

AND2X2 _15251_ (
    .A(_4208__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_4209_)
);

FILL FILL380000x153140 (
);

FILL FILL225720x266760 (
);

FILL FILL331360x340860 (
);

FILL FILL_1__17598_ (
);

AND2X2 _16876_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_5809_)
);

OR2X2 _16456_ (
    .A(_5391_),
    .B(_5394_),
    .Y(_5395_)
);

AND2X2 _16036_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_4982_)
);

AND2X2 _11591_ (
    .A(_1612_),
    .B(_1611_),
    .Y(_1587_[12])
);

AND2X2 _11171_ (
    .A(_1392_),
    .B(_1391_),
    .Y(_1389_[1])
);

FILL FILL_0__17952_ (
);

FILL FILL_0__17532_ (
);

FILL FILL_0__17112_ (
);

FILL FILL114760x69160 (
);

AND2X2 _8798_ (
    .A(_190_),
    .B(_189_),
    .Y(_135_[27])
);

FILL FILL274360x291460 (
);

FILL FILL53200x74100 (
);

NOR2X1 _12796_ (
    .A(_2356_),
    .B(_2360_),
    .Y(_2361_)
);

OR2X2 _12376_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_2048__bF$buf4),
    .Y(_2016_)
);

FILL FILL_0__18737_ (
);

FILL FILL_0__18317_ (
);

AND2X2 _18602_ (
    .A(_6315__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_7509_)
);

FILL FILL_0__13452_ (
);

FILL FILL_0__13032_ (
);

FILL FILL_0__8418_ (
);

FILL FILL196840x74100 (
);

OR2X2 _14942_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [19]),
    .Y(_3974_)
);

FILL FILL_0__14657_ (
);

OR2X2 _14522_ (
    .A(IRWrite_bF$buf3),
    .B(\datapath_1.PCJump [10]),
    .Y(_3754_)
);

OR2X2 _14102_ (
    .A(_3505_),
    .B(_3506_),
    .Y(_3507_)
);

FILL FILL117800x375440 (
);

FILL FILL162640x158080 (
);

FILL FILL_0__18490_ (
);

FILL FILL_0__18070_ (
);

FILL FILL_1__16449_ (
);

OR2X2 _15727_ (
    .A(_4677_),
    .B(_4674_),
    .Y(_4678_)
);

AND2X2 _15307_ (
    .A(_4158__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_4264_)
);

FILL FILL_0__8591_ (
);

AND2X2 _10862_ (
    .A(_1246_),
    .B(_1245_),
    .Y(_1191_[27])
);

FILL FILL_0__10157_ (
);

AND2X2 _10442_ (
    .A(_1026_),
    .B(_1025_),
    .Y(_993_[16])
);

AND2X2 _10022_ (
    .A(_806_),
    .B(_805_),
    .Y(_795_[5])
);

AND2X2 _18199_ (
    .A(_6328__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_7112_)
);

FILL FILL424080x108680 (
);

OR2X2 _19140_ (
    .A(_8037_),
    .B(_8038_),
    .Y(_8039_)
);

FILL FILL227240x370500 (
);

FILL FILL_1__12789_ (
);

FILL FILL504640x83980 (
);

FILL FILL441560x118560 (
);

FILL FILL_0__9796_ (
);

FILL FILL_0__9376_ (
);

OR2X2 _11647_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .B(_1652__bF$buf3),
    .Y(_1650_)
);

OR2X2 _11227_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_1454__bF$buf3),
    .Y(_1430_)
);

FILL FILL_0__12723_ (
);

FILL FILL166440x266760 (
);

OR2X2 _15480_ (
    .A(_4419_),
    .B(_4434_),
    .Y(_4435_)
);

FILL FILL_0__15195_ (
);

NOR2X1 _15060_ (
    .A(_4023_),
    .B(\datapath_1.a3 [4]),
    .Y(_4049_)
);

FILL FILL272080x340860 (
);

FILL FILL_1__14935_ (
);

FILL FILL_0__13928_ (
);

FILL FILL_0__13508_ (
);

AND2X2 _16685_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_5621_)
);

OR2X2 _16265_ (
    .A(_5199_),
    .B(_5206_),
    .Y(_5207_)
);

FILL FILL_0__17341_ (
);

FILL FILL_1__10435_ (
);

DFFSR _12185_ (
    .CLK(clk_bF$buf9),
    .D(_1851_[20]),
    .Q(\datapath_1.regfile_1.regOut[29] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

FILL FILL_1__19133_ (
);

FILL FILL_0__18966_ (
);

FILL FILL16720x321100 (
);

OR2X2 _18831_ (
    .A(_7734_),
    .B(_7733_),
    .Y(_7735_)
);

FILL FILL_0__18546_ (
);

OR2X2 _18411_ (
    .A(_7319_),
    .B(_7320_),
    .Y(_7321_)
);

FILL FILL224960x64220 (
);

FILL FILL_0__13681_ (
);

FILL FILL_0__13261_ (
);

OR2X2 _10918_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .B(_1322__bF$buf2),
    .Y(_1264_)
);

FILL FILL_1__9290_ (
);

FILL FILL164920x222300 (
);

FILL FILL234080x123500 (
);

FILL FILL_1__15053_ (
);

FILL FILL420280x138320 (
);

FILL FILL_0__14886_ (
);

DFFSR _14751_ (
    .CLK(clk_bF$buf94),
    .D(_3804_[28]),
    .Q(\datapath_1.a [28]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL_0__14046_ (
);

OR2X2 _14331_ (
    .A(\datapath_1.ALUResult [30]),
    .B(_3671__bF$buf4),
    .Y(_3667_)
);

FILL FILL163400x34580 (
);

AND2X2 _15956_ (
    .A(_4197__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_4903_)
);

FILL FILL228760x64220 (
);

AND2X2 _15536_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_4490_)
);

OAI21X1 _15116_ (
    .A(_4038_),
    .B(_4094_),
    .C(_4017_),
    .Y(_4095_)
);

OR2X2 _10671_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_1139_)
);

DFFSR _10251_ (
    .CLK(clk_bF$buf28),
    .D(_861_[21]),
    .Q(\datapath_1.regfile_1.regOut[14] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

FILL FILL_0__16612_ (
);

FILL FILL76760x281580 (
);

FILL FILL_0__19084_ (
);

AND2X2 _11876_ (
    .A(_1762_),
    .B(_1761_),
    .Y(_1719_[21])
);

AND2X2 _11456_ (
    .A(_1542_),
    .B(_1541_),
    .Y(_1521_[10])
);

OR2X2 _11036_ (
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .Y(_1387_)
);

FILL FILL_0__17817_ (
);

FILL FILL_0__12952_ (
);

DFFSR _9604_ (
    .CLK(clk_bF$buf60),
    .D(_531_[19]),
    .Q(\datapath_1.regfile_1.regOut[9] [19]),
    .R(rst_bF$buf41),
    .S(vdd)
);

FILL FILL_1__8981_ (
);

FILL FILL_1__14324_ (
);

FILL FILL_0__13317_ (
);

AND2X2 _13602_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3096_)
);

FILL FILL_0_BUFX2_insert1180 (
);

FILL FILL_0_BUFX2_insert1182 (
);

OR2X2 _16494_ (
    .A(_5432_),
    .B(_5431_),
    .Y(_5433_)
);

AND2X2 _16074_ (
    .A(_4195__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_5019_)
);

FILL FILL_0_BUFX2_insert1184 (
);

FILL FILL_0_BUFX2_insert1185 (
);

FILL FILL_0_BUFX2_insert1186 (
);

FILL FILL_0_BUFX2_insert1187 (
);

FILL FILL_0_BUFX2_insert1188 (
);

FILL FILL_0_BUFX2_insert1189 (
);

FILL FILL25840x118560 (
);

FILL FILL_0__17990_ (
);

FILL FILL128440x276640 (
);

FILL FILL_0__17570_ (
);

FILL FILL_1__15949_ (
);

OR2X2 _14807_ (
    .A(vdd),
    .B(_2_[17]),
    .Y(_3904_)
);

FILL FILL435480x103740 (
);

FILL FILL373160x44460 (
);

OR2X2 _17699_ (
    .A(_6612_),
    .B(_6619_),
    .Y(_6620_)
);

AND2X2 _17279_ (
    .A(_6203_),
    .B(_6204_),
    .Y(_6205_)
);

FILL FILL_1__19362_ (
);

FILL FILL125400x64220 (
);

OR2X2 _18640_ (
    .A(_7543_),
    .B(_7546_),
    .Y(_7547_)
);

FILL FILL_0__18355_ (
);

AND2X2 _18220_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_7133_)
);

FILL FILL196840x103740 (
);

FILL FILL_0__13070_ (
);

FILL FILL_1__11869_ (
);

FILL FILL440040x83980 (
);

FILL FILL297160x311220 (
);

AND2X2 _10727_ (
    .A(_1176_),
    .B(_1175_),
    .Y(_1125_[25])
);

AND2X2 _10307_ (
    .A(_956_),
    .B(_955_),
    .Y(_927_[14])
);

FILL FILL190760x256880 (
);

AND2X2 _13199_ (
    .A(_2747_),
    .B(_2742_),
    .Y(_2748_)
);

AND2X2 _19425_ (
    .A(_8319_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.rd1 [31])
);

AND2X2 _19005_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_7906_)
);

FILL FILL_0__14695_ (
);

AND2X2 _14980_ (
    .A(_3999_),
    .B(_3998_),
    .Y(_3936_[31])
);

FILL FILL_0__14275_ (
);

AND2X2 _14560_ (
    .A(_3779_),
    .B(_3778_),
    .Y(_3738_[20])
);

OR2X2 _14140_ (
    .A(_3539_),
    .B(_3538_),
    .Y(_3540_)
);

FILL FILL386840x360620 (
);

FILL FILL_1__16067_ (
);

FILL FILL129200x64220 (
);

FILL FILL211280x0 (
);

AND2X2 _15765_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_4715_)
);

AND2X2 _15345_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [1]),
    .Y(_4302_)
);

FILL FILL_0__10195_ (
);

OR2X2 _10480_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .B(_1058__bF$buf2),
    .Y(_1052_)
);

FILL FILL313120x251940 (
);

OR2X2 _10060_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_860__bF$buf0),
    .Y(_832_)
);

FILL FILL_0__16841_ (
);

FILL FILL_0__16421_ (
);

FILL FILL_0__16001_ (
);

OR2X2 _11685_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_1655_)
);

FILL FILL_1__18213_ (
);

DFFSR _11265_ (
    .CLK(clk_bF$buf44),
    .D(_1389_[3]),
    .Q(\datapath_1.regfile_1.regOut[22] [3]),
    .R(rst_bF$buf16),
    .S(vdd)
);

OR2X2 _17911_ (
    .A(_6821_),
    .B(_6828_),
    .Y(_6829_)
);

FILL FILL_0__17206_ (
);

FILL FILL123120x88920 (
);

FILL FILL85880x9880 (
);

FILL FILL_0__12761_ (
);

FILL FILL505400x98800 (
);

FILL FILL357200x14820 (
);

FILL FILL283480x158080 (
);

AND2X2 _9833_ (
    .A(_720_),
    .B(_719_),
    .Y(_663_[28])
);

AND2X2 _9413_ (
    .A(_500_),
    .B(_499_),
    .Y(_465_[17])
);

FILL FILL_1__8790_ (
);

FILL FILL169480x182780 (
);

FILL FILL335160x74100 (
);

FILL FILL21280x375440 (
);

FILL FILL267520x49400 (
);

FILL FILL_0__13546_ (
);

OR2X2 _13831_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [5]),
    .Y(_3287_)
);

FILL FILL_0__13126_ (
);

OR2X2 _13411_ (
    .A(_2387__bF$buf0),
    .B(_2946_),
    .Y(_2947_)
);

FILL FILL431680x0 (
);

FILL FILL224200x202540 (
);

DFFSR _14616_ (
    .CLK(clk_bF$buf2),
    .D(_3738_[22]),
    .Q(\datapath_1.PCJump [24]),
    .R(rst_bF$buf33),
    .S(vdd)
);

FILL FILL410400x217360 (
);

OR2X2 _17088_ (
    .A(_6015_),
    .B(_6016_),
    .Y(_6017_)
);

FILL FILL167200x153140 (
);

FILL FILL_0__18584_ (
);

FILL FILL_0__18164_ (
);

OR2X2 _10956_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_1289_)
);

OR2X2 _10536_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_1069_)
);

DFFSR _10116_ (
    .CLK(clk_bF$buf89),
    .D(_795_[15]),
    .Q(\datapath_1.regfile_1.regOut[13] [15]),
    .R(rst_bF$buf24),
    .S(vdd)
);

FILL FILL_0__11612_ (
);

FILL FILL_1__15091_ (
);

FILL FILL_0__19369_ (
);

AND2X2 _19234_ (
    .A(_6250__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_8131_)
);

FILL FILL_0__14084_ (
);

FILL FILL72200x207480 (
);

FILL FILL_0__12817_ (
);

FILL FILL376200x118560 (
);

AND2X2 _15994_ (
    .A(_4940_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [11])
);

FILL FILL_0__15289_ (
);

OR2X2 _15574_ (
    .A(_4525_),
    .B(_4526_),
    .Y(_4527_)
);

AND2X2 _15154_ (
    .A(_4118_),
    .B(_4117_),
    .Y(\datapath_1.regfile_1.regEn [25])
);

FILL FILL_0__16650_ (
);

AND2X2 _16779_ (
    .A(_4172__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [24]),
    .Y(_5713_)
);

OR2X2 _16359_ (
    .A(_5299_),
    .B(_5296_),
    .Y(_5300_)
);

FILL FILL_1__18862_ (
);

OR2X2 _11494_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .B(_1586__bF$buf3),
    .Y(_1568_)
);

OR2X2 _11074_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_1388__bF$buf0),
    .Y(_1348_)
);

FILL FILL_0__17435_ (
);

AND2X2 _17720_ (
    .A(_6289__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_6641_)
);

AND2X2 _17300_ (
    .A(_6225_),
    .B(\datapath_1.PCJump [24]),
    .Y(_6226_)
);

FILL FILL_0__12570_ (
);

FILL FILL_0__12150_ (
);

FILL FILL370880x256880 (
);

FILL FILL_1__10529_ (
);

OR2X2 _9642_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_613_)
);

DFFSR _9222_ (
    .CLK(clk_bF$buf35),
    .D(_333_[24]),
    .Q(\datapath_1.regfile_1.regOut[6] [24]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL110960x128440 (
);

AND2X2 _12699_ (
    .A(_2262_),
    .B(_2263_),
    .Y(_2264_)
);

FILL FILL_1__19227_ (
);

OR2X2 _12279_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_1971_)
);

FILL FILL_1__14782_ (
);

OR2X2 _18925_ (
    .A(_7823_),
    .B(_7826_),
    .Y(_7827_)
);

AND2X2 _18505_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_7414_)
);

FILL FILL_0__13775_ (
);

AND2X2 _13640_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[7]),
    .Y(_3128_)
);

OR2X2 _13220_ (
    .A(_2387__bF$buf3),
    .B(_2766_),
    .Y(_2767_)
);

FILL FILL104880x14820 (
);

FILL FILL432440x281580 (
);

FILL FILL107920x79040 (
);

FILL FILL124640x29640 (
);

FILL FILL_1__15567_ (
);

AND2X2 _14845_ (
    .A(_3929_),
    .B(_3928_),
    .Y(_3870_[29])
);

AND2X2 _14425_ (
    .A(_3709_),
    .B(_3708_),
    .Y(_3672_[18])
);

AND2X2 _14005_ (
    .A(_3350__bF$buf3),
    .B(_2_[12]),
    .Y(_3424_)
);

FILL FILL_0__15501_ (
);

FILL FILL_0__18393_ (
);

FILL FILL391400x311220 (
);

FILL FILL_0__8494_ (
);

DFFSR _10765_ (
    .CLK(clk_bF$buf16),
    .D(_1125_[19]),
    .Q(\datapath_1.regfile_1.regOut[18] [19]),
    .R(rst_bF$buf20),
    .S(vdd)
);

FILL FILL_1__17713_ (
);

OR2X2 _10345_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .B(_992__bF$buf4),
    .Y(_982_)
);

FILL FILL_0__16706_ (
);

FILL FILL313880x197600 (
);

FILL FILL_0__11841_ (
);

FILL FILL_0__11001_ (
);

FILL FILL_0__19178_ (
);

OR2X2 _19463_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_8344_)
);

AND2X2 _19043_ (
    .A(_6259__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_7943_)
);

FILL FILL128440x29640 (
);

OR2X2 _8913_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_247_)
);

FILL FILL_1_BUFX2_insert411 (
);

INVX1 _12911_ (
    .A(_2330_),
    .Y(_2476_)
);

FILL FILL_0__12626_ (
);

FILL FILL_0__12206_ (
);

FILL FILL_1_BUFX2_insert419 (
);

FILL FILL232560x44460 (
);

FILL FILL_0__15098_ (
);

OR2X2 _15383_ (
    .A(_4335_),
    .B(_4338_),
    .Y(_4339_)
);

FILL FILL43320x242060 (
);

FILL FILL115520x83980 (
);

OR2X2 _16588_ (
    .A(_5523_),
    .B(_5524_),
    .Y(_5525_)
);

OR2X2 _16168_ (
    .A(_5104_),
    .B(_5111_),
    .Y(_5112_)
);

FILL FILL_0__17664_ (
);

DFFSR _9871_ (
    .CLK(clk_bF$buf61),
    .D(_663_[28]),
    .Q(\datapath_1.regfile_1.regOut[11] [28]),
    .R(rst_bF$buf58),
    .S(vdd)
);

OR2X2 _9451_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .B(_530__bF$buf1),
    .Y(_526_)
);

OR2X2 _9031_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .B(_332__bF$buf0),
    .Y(_306_)
);

OR2X2 _12088_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_1916__bF$buf2),
    .Y(_1864_)
);

FILL FILL370880x29640 (
);

FILL FILL_0__18869_ (
);

OR2X2 _18734_ (
    .A(_7637_),
    .B(_7638_),
    .Y(_7639_)
);

OR2X2 _18314_ (
    .A(_7224_),
    .B(_7225_),
    .Y(_7226_)
);

FILL FILL_0__18029_ (
);

FILL FILL_0__13164_ (
);

FILL FILL47120x29640 (
);

FILL FILL_1__9193_ (
);

FILL FILL_0__9911_ (
);

FILL FILL482600x247000 (
);

AND2X2 _19519_ (
    .A(_8381_),
    .B(_8380_),
    .Y(_8320_[30])
);

FILL FILL_0__14789_ (
);

OR2X2 _14654_ (
    .A(vdd),
    .B(\datapath_1.a [9]),
    .Y(_3822_)
);

FILL FILL104120x128440 (
);

OR2X2 _14234_ (
    .A(\datapath_1.Data [30]),
    .B(_3605__bF$buf3),
    .Y(_3601_)
);

FILL FILL378480x217360 (
);

FILL FILL140600x301340 (
);

FILL FILL_0__15730_ (
);

FILL FILL_0__15310_ (
);

FILL FILL91960x316160 (
);

FILL FILL199120x172900 (
);

FILL FILL_1__11296_ (
);

AND2X2 _15859_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_4808_)
);

OR2X2 _15439_ (
    .A(_4392_),
    .B(_4393_),
    .Y(_4394_)
);

OAI21X1 _15019_ (
    .A(_4004_),
    .B(_4007_),
    .C(\datapath_1.a3 [4]),
    .Y(_4008_)
);

FILL FILL150480x83980 (
);

AND2X2 _10994_ (
    .A(_1314_),
    .B(_1313_),
    .Y(_1257_[28])
);

FILL FILL_0__10289_ (
);

AND2X2 _10574_ (
    .A(_1094_),
    .B(_1093_),
    .Y(_1059_[17])
);

AND2X2 _10154_ (
    .A(_874_),
    .B(_873_),
    .Y(_861_[6])
);

FILL FILL462080x69160 (
);

FILL FILL_0__16935_ (
);

FILL FILL_0__16515_ (
);

OR2X2 _16800_ (
    .A(_5730_),
    .B(_5733_),
    .Y(_5734_)
);

FILL FILL_0__11230_ (
);

FILL FILL325280x93860 (
);

AND2X2 _19272_ (
    .A(_6287__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_8169_)
);

FILL FILL170240x163020 (
);

OR2X2 _8722_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .B(_200__bF$buf3),
    .Y(_140_)
);

FILL FILL135280x326040 (
);

FILL FILL22040x128440 (
);

FILL FILL_1__18727_ (
);

DFFSR _11779_ (
    .CLK(clk_bF$buf16),
    .D(_1653_[1]),
    .Q(\datapath_1.regfile_1.regOut[26] [1]),
    .R(rst_bF$buf20),
    .S(vdd)
);

OR2X2 _11359_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .B(_1520__bF$buf1),
    .Y(_1498_)
);

FILL FILL430920x330980 (
);

FILL FILL_1__13442_ (
);

NAND3X1 _12720_ (
    .A(_2281_),
    .B(_2277_),
    .C(_2284_),
    .Y(_2285_)
);

FILL FILL_0__12015_ (
);

DFFSR _12300_ (
    .CLK(clk_bF$buf7),
    .D(_1917_[6]),
    .Q(\datapath_1.regfile_1.regOut[30] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

NAND2X1 _15192_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_4150_)
);

FILL FILL489440x69160 (
);

FILL FILL422560x24700 (
);

OR2X2 _9927_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_763_)
);

OR2X2 _9507_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_543_)
);

FILL FILL_1__8884_ (
);

FILL FILL65360x79040 (
);

FILL FILL292600x217360 (
);

AND2X2 _13925_ (
    .A(_3344__bF$buf2),
    .B(gnd),
    .Y(_3355_)
);

OR2X2 _13505_ (
    .A(ALUOut[5]),
    .B(_3079__bF$buf0),
    .Y(_3025_)
);

AND2X2 _16397_ (
    .A(_4160__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_5337_)
);

FILL FILL_1__18480_ (
);

FILL FILL_1__9249_ (
);

FILL FILL_0__17473_ (
);

FILL FILL_0__17053_ (
);

FILL FILL_1__10567_ (
);

FILL FILL186960x355680 (
);

AND2X2 _9680_ (
    .A(_638_),
    .B(_637_),
    .Y(_597_[20])
);

AND2X2 _9260_ (
    .A(_418_),
    .B(_417_),
    .Y(_399_[9])
);

FILL FILL_1_CLKBUF1_insert125 (
);

FILL FILL_1_CLKBUF1_insert127 (
);

FILL FILL_1_CLKBUF1_insert129 (
);

FILL FILL_0__10921_ (
);

FILL FILL14440x143260 (
);

FILL FILL_0__18678_ (
);

AND2X2 _18963_ (
    .A(_6211__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_7865_)
);

OR2X2 _18543_ (
    .A(_7450_),
    .B(_7447_),
    .Y(_7451_)
);

FILL FILL_0__18258_ (
);

OR2X2 _18123_ (
    .A(_7006_),
    .B(_7037_),
    .Y(_7038_)
);

FILL FILL_0__13393_ (
);

FILL FILL130720x256880 (
);

FILL FILL_0__11706_ (
);

FILL FILL_0__9300_ (
);

FILL FILL_1__15185_ (
);

AND2X2 _19328_ (
    .A(_6287__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_8224_)
);

DFFSR _14883_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[31]),
    .Q(_2_[31]),
    .R(rst_bF$buf61),
    .S(vdd)
);

OR2X2 _14463_ (
    .A(memoryOutData[31]),
    .B(_3737__bF$buf1),
    .Y(_3735_)
);

OR2X2 _14043_ (
    .A(_3456_),
    .B(_3453_),
    .Y(\datapath_1.alu_1.ALUInB [17])
);

FILL FILL335160x291460 (
);

FILL FILL_1__13918_ (
);

FILL FILL427120x247000 (
);

AND2X2 _15668_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_4620_)
);

FILL FILL433200x93860 (
);

OR2X2 _15248_ (
    .A(_4205_),
    .B(_4199_),
    .Y(_4206_)
);

FILL FILL54720x103740 (
);

FILL FILL_0__10098_ (
);

FILL FILL_1__17331_ (
);

DFFSR _10383_ (
    .CLK(clk_bF$buf97),
    .D(_927_[24]),
    .Q(\datapath_1.regfile_1.regOut[15] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

OR2X2 _19081_ (
    .A(_7980_),
    .B(_7973_),
    .Y(_7981_)
);

DFFSR _8951_ (
    .CLK(clk_bF$buf71),
    .D(_201_[11]),
    .Q(\datapath_1.regfile_1.regOut[4] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

AND2X2 _8531_ (
    .A(_52_),
    .B(_51_),
    .Y(_3_[24])
);

AND2X2 _11588_ (
    .A(_1610_),
    .B(_1609_),
    .Y(_1587_[11])
);

AND2X2 _11168_ (
    .A(_1390_),
    .B(_1453_),
    .Y(_1389_[0])
);

FILL FILL71440x340860 (
);

FILL FILL_1__13671_ (
);

FILL FILL_0__17949_ (
);

FILL FILL_0__17529_ (
);

OR2X2 _17814_ (
    .A(_6731_),
    .B(_6732_),
    .Y(_6733_)
);

FILL FILL_0__12664_ (
);

DFFSR _9736_ (
    .CLK(clk_bF$buf72),
    .D(_597_[22]),
    .Q(\datapath_1.regfile_1.regOut[10] [22]),
    .R(rst_bF$buf2),
    .S(vdd)
);

OR2X2 _9316_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .B(_464__bF$buf4),
    .Y(_456_)
);

FILL FILL109440x182780 (
);

FILL FILL66880x138320 (
);

FILL FILL493240x148200 (
);

FILL FILL_0__13869_ (
);

AND2X2 _13734_ (
    .A(_3087__bF$buf2),
    .B(\datapath_1.ALUResult [20]),
    .Y(_3209_)
);

AND2X2 _13314_ (
    .A(_2854_),
    .B(_2852_),
    .Y(_2855_)
);

FILL FILL_0__13029_ (
);

FILL FILL415720x207480 (
);

FILL FILL_0__14810_ (
);

FILL FILL6840x9880 (
);

FILL FILL_0__17282_ (
);

FILL FILL153520x74100 (
);

FILL FILL132240x360620 (
);

OR2X2 _14939_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [18]),
    .Y(_3972_)
);

OR2X2 _14519_ (
    .A(IRWrite_bF$buf3),
    .B(\datapath_1.PCJump [9]),
    .Y(_3752_)
);

FILL FILL_0__10730_ (
);

OR2X2 _18772_ (
    .A(_7661_),
    .B(_7676_),
    .Y(_7677_)
);

FILL FILL_0__18487_ (
);

AND2X2 _18352_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [15]),
    .Y(_7263_)
);

FILL FILL481840x242060 (
);

FILL FILL44840x192660 (
);

FILL FILL_1__17807_ (
);

AND2X2 _10859_ (
    .A(_1244_),
    .B(_1243_),
    .Y(_1191_[26])
);

AND2X2 _10439_ (
    .A(_1024_),
    .B(_1023_),
    .Y(_993_[15])
);

FILL FILL286520x202540 (
);

AND2X2 _10019_ (
    .A(_804_),
    .B(_803_),
    .Y(_795_[4])
);

FILL FILL364800x74100 (
);

FILL FILL436240x365560 (
);

DFFSR _11800_ (
    .CLK(clk_bF$buf26),
    .D(_1653_[22]),
    .Q(\datapath_1.regfile_1.regOut[26] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL267520x360620 (
);

AND2X2 _19557_ (
    .A(Branch),
    .B(ALUZero),
    .Y(_8388_)
);

OR2X2 _19137_ (
    .A(_8035_),
    .B(_8032_),
    .Y(_8036_)
);

AND2X2 _14692_ (
    .A(_3847_),
    .B(_3846_),
    .Y(_3804_[21])
);

AND2X2 _14272_ (
    .A(_3627_),
    .B(_3626_),
    .Y(_3606_[10])
);

FILL FILL50160x360620 (
);

FILL FILL258400x335920 (
);

FILL FILL_1__13307_ (
);

FILL FILL158840x9880 (
);

OR2X2 _15897_ (
    .A(_4829_),
    .B(_4844_),
    .Y(_4845_)
);

OR2X2 _15477_ (
    .A(_4430_),
    .B(_4431_),
    .Y(_4432_)
);

AND2X2 _15057_ (
    .A(_4044_),
    .B(_4045_),
    .Y(_4046_)
);

FILL FILL_1__17980_ (
);

OR2X2 _10192_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .B(_926__bF$buf0),
    .Y(_900_)
);

FILL FILL_0__16553_ (
);

FILL FILL_0__16133_ (
);

OR2X2 _8760_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_165_)
);

DFFSR _11397_ (
    .CLK(clk_bF$buf7),
    .D(_1455_[6]),
    .Q(\datapath_1.regfile_1.regOut[23] [6]),
    .R(rst_bF$buf48),
    .S(vdd)
);

FILL FILL411920x237120 (
);

FILL FILL_1__13060_ (
);

FILL FILL_0__17758_ (
);

AND2X2 _17623_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_6545_)
);

FILL FILL_0__17338_ (
);

AND2X2 _17203_ (
    .A(_4214__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_6131_)
);

FILL FILL_0__12893_ (
);

FILL FILL_0__12473_ (
);

FILL FILL316160x330980 (
);

AND2X2 _9965_ (
    .A(_788_),
    .B(_787_),
    .Y(_729_[29])
);

AND2X2 _9545_ (
    .A(_568_),
    .B(_567_),
    .Y(_531_[18])
);

AND2X2 _9125_ (
    .A(_348_),
    .B(_347_),
    .Y(_333_[7])
);

FILL FILL333640x340860 (
);

FILL FILL178600x98800 (
);

FILL FILL_0__8800_ (
);

FILL FILL_1__14685_ (
);

OR2X2 _18828_ (
    .A(_7731_),
    .B(_7728_),
    .Y(_7732_)
);

FILL FILL_0_BUFX2_insert450 (
);

FILL FILL_0_BUFX2_insert451 (
);

OR2X2 _18408_ (
    .A(_7317_),
    .B(_7316_),
    .Y(_7318_)
);

FILL FILL_0_BUFX2_insert452 (
);

FILL FILL_0_BUFX2_insert453 (
);

FILL FILL_0_BUFX2_insert454 (
);

AND2X2 _13963_ (
    .A(_3350__bF$buf3),
    .B(_2_[6]),
    .Y(_3388_)
);

FILL FILL_0__13678_ (
);

FILL FILL_0__13258_ (
);

OR2X2 _13543_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [18]),
    .Y(_3050_)
);

NAND2X1 _13123_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2676_)
);

FILL FILL_0_BUFX2_insert456 (
);

FILL FILL_0_BUFX2_insert458 (
);

FILL FILL192280x74100 (
);

FILL FILL276640x291460 (
);

FILL FILL_0__17091_ (
);

DFFSR _14748_ (
    .CLK(clk_bF$buf58),
    .D(_3804_[25]),
    .Q(\datapath_1.a [25]),
    .R(rst_bF$buf15),
    .S(vdd)
);

OR2X2 _14328_ (
    .A(\datapath_1.ALUResult [29]),
    .B(_3671__bF$buf3),
    .Y(_3665_)
);

FILL FILL_1__16831_ (
);

FILL FILL377720x138320 (
);

FILL FILL_0__15824_ (
);

FILL FILL_0__15404_ (
);

AND2X2 _18581_ (
    .A(_6244__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_7488_)
);

OR2X2 _18161_ (
    .A(_7074_),
    .B(_7073_),
    .Y(_7075_)
);

FILL FILL_0_CLKBUF1_insert1170 (
);

FILL FILL_0_CLKBUF1_insert1172 (
);

FILL FILL_0_CLKBUF1_insert1173 (
);

FILL FILL_0_CLKBUF1_insert1174 (
);

FILL FILL_0_CLKBUF1_insert1175 (
);

FILL FILL_0_CLKBUF1_insert1176 (
);

FILL FILL_0_CLKBUF1_insert1178 (
);

FILL FILL221920x207480 (
);

OR2X2 _10668_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_1137_)
);

DFFSR _10248_ (
    .CLK(clk_bF$buf106),
    .D(_861_[18]),
    .Q(\datapath_1.regfile_1.regOut[14] [18]),
    .R(rst_bF$buf0),
    .S(vdd)
);

FILL FILL122360x103740 (
);

FILL FILL_0__11744_ (
);

FILL FILL199120x335920 (
);

OR2X2 _19366_ (
    .A(_8259_),
    .B(_8260_),
    .Y(_8261_)
);

OR2X2 _14081_ (
    .A(_3487_),
    .B(_3488_),
    .Y(_3489_)
);

DFFSR _8816_ (
    .CLK(clk_bF$buf104),
    .D(_135_[5]),
    .Q(\datapath_1.regfile_1.regOut[3] [5]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL481080x286520 (
);

FILL FILL_1__13956_ (
);

FILL FILL_1__13536_ (
);

FILL FILL398240x296400 (
);

FILL FILL48640x232180 (
);

NOR2X1 _12814_ (
    .A(_2375_),
    .B(_2378_),
    .Y(_2379_)
);

FILL FILL_0__12529_ (
);

FILL FILL_0__12109_ (
);

FILL FILL38000x192660 (
);

OR2X2 _15286_ (
    .A(_4238_),
    .B(_4243_),
    .Y(_4244_)
);

FILL FILL39520x207480 (
);

FILL FILL426360x108680 (
);

FILL FILL_0__16782_ (
);

FILL FILL_1__18154_ (
);

FILL FILL168720x266760 (
);

FILL FILL_0__17987_ (
);

OR2X2 _17852_ (
    .A(_6769_),
    .B(_6770_),
    .Y(_6771_)
);

AND2X2 _17432_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_6357_)
);

FILL FILL_0__17147_ (
);

AND2X2 _17012_ (
    .A(_4208__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_5943_)
);

FILL FILL_0__12282_ (
);

FILL FILL92720x59280 (
);

OR2X2 _9774_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_681_)
);

DFFSR _9354_ (
    .CLK(clk_bF$buf36),
    .D(_399_[27]),
    .Q(\datapath_1.regfile_1.regOut[7] [27]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL505400x143260 (
);

AND2X2 _18637_ (
    .A(_6323__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_7544_)
);

OR2X2 _18217_ (
    .A(_7126_),
    .B(_7129_),
    .Y(_7130_)
);

FILL FILL_0__13487_ (
);

OR2X2 _13772_ (
    .A(_3241_),
    .B(_3238_),
    .Y(\datapath_1.mux_pcsrc.dout [25])
);

XOR2X1 _13352_ (
    .A(_2196_),
    .B(_2890_),
    .Y(_2891_)
);

FILL FILL_0__13067_ (
);

FILL FILL291080x256880 (
);

FILL FILL437000x29640 (
);

FILL FILL_0__9814_ (
);

FILL FILL401280x207480 (
);

AND2X2 _14977_ (
    .A(_3997_),
    .B(_3996_),
    .Y(_3936_[30])
);

AND2X2 _14557_ (
    .A(_3777_),
    .B(_3776_),
    .Y(_3738_[19])
);

OR2X2 _14137_ (
    .A(_3535_),
    .B(_3536_),
    .Y(_3537_)
);

FILL FILL_0__15633_ (
);

FILL FILL490960x177840 (
);

AND2X2 _18390_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_7300_)
);

FILL FILL266000x19760 (
);

FILL FILL441560x301340 (
);

DFFSR _10897_ (
    .CLK(clk_bF$buf26),
    .D(_1191_[22]),
    .Q(\datapath_1.regfile_1.regOut[19] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL_1__17845_ (
);

OR2X2 _10477_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_1058__bF$buf1),
    .Y(_1050_)
);

OR2X2 _10057_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_860__bF$buf4),
    .Y(_830_)
);

FILL FILL_1__12140_ (
);

FILL FILL_0__16418_ (
);

AND2X2 _16703_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_5638_)
);

FILL FILL_0__11973_ (
);

FILL FILL_0__11553_ (
);

FILL FILL221920x345800 (
);

OR2X2 _19175_ (
    .A(_8071_),
    .B(_8072_),
    .Y(_8073_)
);

FILL FILL403560x296400 (
);

FILL FILL370120x34580 (
);

OR2X2 _8625_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_95_)
);

FILL FILL253080x360620 (
);

AND2X2 _17908_ (
    .A(_6297__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_6826_)
);

FILL FILL268280x14820 (
);

FILL FILL_0__12758_ (
);

NAND2X1 _12623_ (
    .A(_2186_),
    .B(_2187_),
    .Y(_2188_)
);

FILL FILL_0__12338_ (
);

AND2X2 _12203_ (
    .A(_1920_),
    .B(_1919_),
    .Y(_1917_[1])
);

FILL FILL80560x207480 (
);

AND2X2 _15095_ (
    .A(_4078_),
    .B(_4029_),
    .Y(\datapath_1.regfile_1.regEn [6])
);

FILL FILL143640x93860 (
);

FILL FILL_0__16591_ (
);

FILL FILL_0__16171_ (
);

FILL FILL133000x113620 (
);

OR2X2 _13828_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [4]),
    .Y(_3285_)
);

AND2X2 _13408_ (
    .A(_2942_),
    .B(_2943_),
    .Y(_2944_)
);

FILL FILL_0__14904_ (
);

FILL FILL_0__17796_ (
);

OR2X2 _17661_ (
    .A(_6581_),
    .B(_6582_),
    .Y(_6583_)
);

FILL FILL_0__17376_ (
);

OR2X2 _17241_ (
    .A(_6152_),
    .B(_6167_),
    .Y(_6168_)
);

FILL FILL_0__12091_ (
);

OR2X2 _9583_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .B(_596__bF$buf1),
    .Y(_594_)
);

OR2X2 _9163_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_398__bF$buf1),
    .Y(_374_)
);

FILL FILL_1__11831_ (
);

FILL FILL323000x370500 (
);

FILL FILL_1__19168_ (
);

FILL FILL437000x118560 (
);

OR2X2 _18866_ (
    .A(_7768_),
    .B(_7767_),
    .Y(_7769_)
);

FILL FILL_0_BUFX2_insert830 (
);

FILL FILL_0_BUFX2_insert831 (
);

OR2X2 _18446_ (
    .A(_7348_),
    .B(_7355_),
    .Y(_7356_)
);

FILL FILL_0_BUFX2_insert832 (
);

AND2X2 _18026_ (
    .A(_6272__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_6942_)
);

FILL FILL_0_BUFX2_insert833 (
);

FILL FILL300960x271700 (
);

AND2X2 _13581_ (
    .A(_3075_),
    .B(_3074_),
    .Y(_1_[30])
);

FILL FILL_0_BUFX2_insert835 (
);

OR2X2 _13161_ (
    .A(_2711_),
    .B(_2710_),
    .Y(_2712_)
);

FILL FILL_0_BUFX2_insert837 (
);

FILL FILL_0_BUFX2_insert839 (
);

FILL FILL_0__19102_ (
);

FILL FILL228000x49400 (
);

FILL FILL59280x133380 (
);

FILL FILL_0__9623_ (
);

FILL FILL_0__11609_ (
);

FILL FILL437760x103740 (
);

OR2X2 _14786_ (
    .A(vdd),
    .B(_2_[10]),
    .Y(_3890_)
);

DFFSR _14366_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[30]),
    .Q(ALUOut[30]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL148200x64220 (
);

FILL FILL_0__15022_ (
);

FILL FILL299440x311220 (
);

FILL FILL454480x340860 (
);

FILL FILL82080x311220 (
);

AND2X2 _10286_ (
    .A(_942_),
    .B(_941_),
    .Y(_927_[7])
);

FILL FILL_0__16647_ (
);

AND2X2 _16932_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_5864_)
);

OR2X2 _16512_ (
    .A(_5448_),
    .B(_5449_),
    .Y(_5450_)
);

FILL FILL_0__16227_ (
);

FILL FILL_0__11362_ (
);

OR2X2 _8854_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_266__bF$buf0),
    .Y(_208_)
);

BUFX2 _8434_ (
    .A(_2_[10]),
    .Y(memoryWriteData[10])
);

FILL FILL_1__18019_ (
);

AND2X2 _17717_ (
    .A(_6287__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_6638_)
);

FILL FILL_0__12987_ (
);

FILL FILL120080x247000 (
);

FILL FILL150480x158080 (
);

OR2X2 _12852_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2417_)
);

DFFSR _12432_ (
    .CLK(clk_bF$buf24),
    .D(_1983_[9]),
    .Q(\datapath_1.regfile_1.regOut[31] [9]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_0__12147_ (
);

OR2X2 _12012_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_1833_)
);

OR2X2 _9639_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_611_)
);

DFFSR _9219_ (
    .CLK(clk_bF$buf106),
    .D(_333_[21]),
    .Q(\datapath_1.regfile_1.regOut[6] [21]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL329840x212420 (
);

FILL FILL109440x296400 (
);

AND2X2 _13637_ (
    .A(_3089__bF$buf0),
    .B(gnd),
    .Y(_3126_)
);

NAND2X1 _13217_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2764_)
);

FILL FILL_1__15300_ (
);

AND2X2 _17890_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_6808_)
);

OR2X2 _17470_ (
    .A(_6391_),
    .B(_6394_),
    .Y(_6395_)
);

AND2X2 _17050_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_5980_)
);

FILL FILL55480x163020 (
);

FILL FILL_1__10699_ (
);

FILL FILL177840x123500 (
);

FILL FILL_1__16925_ (
);

AND2X2 _9392_ (
    .A(_486_),
    .B(_485_),
    .Y(_465_[10])
);

FILL FILL_0__15918_ (
);

FILL FILL291080x326040 (
);

OR2X2 _18675_ (
    .A(_7580_),
    .B(_7566_),
    .Y(_7581_)
);

AND2X2 _18255_ (
    .A(_7167_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.rd1 [13])
);

NAND3X1 _13390_ (
    .A(_2383_),
    .B(_2397_),
    .C(_2926_),
    .Y(_2927_)
);

FILL FILL_0__19331_ (
);

FILL FILL158080x187720 (
);

FILL FILL269800x4940 (
);

FILL FILL450680x370500 (
);

FILL FILL_0__11838_ (
);

FILL FILL_0__9432_ (
);

FILL FILL_0__9012_ (
);

OR2X2 _11703_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_1667_)
);

DFFSR _14595_ (
    .CLK(clk_bF$buf65),
    .D(_3738_[1]),
    .Q(\aluControl_1.inst [1]),
    .R(rst_bF$buf91),
    .S(vdd)
);

AND2X2 _14175_ (
    .A(_3561_),
    .B(_3560_),
    .Y(\datapath_1.mux_wd3.dout [10])
);

FILL FILL217360x306280 (
);

FILL FILL288800x4940 (
);

FILL FILL_0__15671_ (
);

FILL FILL_0__15251_ (
);

FILL FILL330600x123500 (
);

FILL FILL234840x316160 (
);

AND2X2 _12908_ (
    .A(_2470_),
    .B(_2472_),
    .Y(_2473_)
);

FILL FILL_1_BUFX2_insert382 (
);

FILL FILL_1_BUFX2_insert384 (
);

FILL FILL_1_BUFX2_insert386 (
);

OR2X2 _10095_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_855_)
);

FILL FILL_0__16876_ (
);

AND2X2 _16741_ (
    .A(_4142__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_5676_)
);

FILL FILL_0__16456_ (
);

OR2X2 _16321_ (
    .A(_5258_),
    .B(_5261_),
    .Y(_5262_)
);

FILL FILL_0__11591_ (
);

AND2X2 _8663_ (
    .A(_120_),
    .B(_119_),
    .Y(_69_[25])
);

FILL FILL9120x153140 (
);

FILL FILL_1__18668_ (
);

FILL FILL_1__18248_ (
);

AND2X2 _17946_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_6863_)
);

AND2X2 _17526_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_6450_)
);

AND2X2 _17106_ (
    .A(_4210__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_6035_)
);

FILL FILL_0__12796_ (
);

OR2X2 _12661_ (
    .A(_2225_),
    .B(_2210_),
    .Y(_2226_)
);

OR2X2 _12241_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_1982__bF$buf2),
    .Y(_1946_)
);

DFFSR _9868_ (
    .CLK(clk_bF$buf93),
    .D(_663_[25]),
    .Q(\datapath_1.regfile_1.regOut[11] [25]),
    .R(rst_bF$buf41),
    .S(vdd)
);

OR2X2 _9448_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .B(_530__bF$buf1),
    .Y(_524_)
);

OR2X2 _9028_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .B(_332__bF$buf1),
    .Y(_304_)
);

AND2X2 _13866_ (
    .A(_3310_),
    .B(_3309_),
    .Y(\datapath_1.alu_1.ALUInA [16])
);

AND2X2 _13446_ (
    .A(_2978_),
    .B(_2763_),
    .Y(_2979_)
);

OR2X2 _13026_ (
    .A(_2584_),
    .B(_2583_),
    .Y(_2585_)
);

FILL FILL_0__14942_ (
);

FILL FILL103360x79040 (
);

FILL FILL_0__9908_ (
);

FILL FILL121600x251940 (
);

FILL FILL_1__16314_ (
);

FILL FILL_0__10862_ (
);

FILL FILL_0__10442_ (
);

FILL FILL_0__18199_ (
);

OR2X2 _18484_ (
    .A(_7391_),
    .B(_7392_),
    .Y(_7393_)
);

INVX1 _18064_ (
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_6979_)
);

FILL FILL378480x59280 (
);

FILL FILL_0__19140_ (
);

FILL FILL_1__12654_ (
);

FILL FILL_0__9661_ (
);

FILL FILL_0__9241_ (
);

DFFSR _11932_ (
    .CLK(clk_bF$buf80),
    .D(_1719_[25]),
    .Q(\datapath_1.regfile_1.regOut[27] [25]),
    .R(rst_bF$buf76),
    .S(vdd)
);

OR2X2 _11512_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .B(_1586__bF$buf4),
    .Y(_1580_)
);

AND2X2 _19269_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_8166_)
);

FILL FILL271320x123500 (
);

OR2X2 _8719_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .B(_200__bF$buf4),
    .Y(_138_)
);

FILL FILL251560x44460 (
);

FILL FILL_0__15060_ (
);

FILL FILL210520x232180 (
);

FILL FILL503880x365560 (
);

FILL FILL338200x296400 (
);

FILL FILL247760x355680 (
);

XNOR2X1 _12717_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2282_)
);

FILL FILL17480x360620 (
);

FILL FILL426360x54340 (
);

FILL FILL_1_BUFX2_insert52 (
);

FILL FILL_1_BUFX2_insert54 (
);

AND2X2 _15189_ (
    .A(_4146__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_4147_)
);

FILL FILL_1_BUFX2_insert56 (
);

FILL FILL_1__17272_ (
);

FILL FILL34960x370500 (
);

AND2X2 _16970_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_5901_)
);

OR2X2 _16550_ (
    .A(_5487_),
    .B(_5486_),
    .Y(_5488_)
);

FILL FILL_0__16265_ (
);

AND2X2 _16130_ (
    .A(_4203__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_5074_)
);

FILL FILL_1__9822_ (
);

OR2X2 _8892_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_233_)
);

FILL FILL114000x247000 (
);

OR2X2 _8472_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_13_)
);

FILL FILL_1__10720_ (
);

FILL FILL110960x311220 (
);

FILL FILL_1__18897_ (
);

OR2X2 _17755_ (
    .A(_6673_),
    .B(_6674_),
    .Y(_6675_)
);

FILL FILL406600x202540 (
);

OR2X2 _17335_ (
    .A(_6260_),
    .B(_6256_),
    .Y(_6261_)
);

FILL FILL255360x44460 (
);

OR2X2 _12890_ (
    .A(_2454_),
    .B(_2452_),
    .Y(_2455_)
);

NOR2X1 _12470_ (
    .A(\aluControl_1.inst [3]),
    .B(\aluControl_1.inst [2]),
    .Y(_2063_)
);

DFFSR _12050_ (
    .CLK(clk_bF$buf85),
    .D(_1785_[14]),
    .Q(\datapath_1.regfile_1.regOut[28] [14]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL_0__18831_ (
);

FILL FILL_0__18411_ (
);

FILL FILL345800x83980 (
);

AND2X2 _9677_ (
    .A(_636_),
    .B(_635_),
    .Y(_597_[19])
);

AND2X2 _9257_ (
    .A(_416_),
    .B(_415_),
    .Y(_399_[8])
);

FILL FILL97280x237120 (
);

FILL FILL_0__8512_ (
);

FILL FILL_1_BUFX2_insert1142 (
);

FILL FILL218120x261820 (
);

FILL FILL_1_BUFX2_insert1144 (
);

AND2X2 _13675_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[12]),
    .Y(_3158_)
);

NAND2X1 _13255_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2800_)
);

FILL FILL_1_BUFX2_insert1146 (
);

FILL FILL404320x276640 (
);

FILL FILL285000x326040 (
);

FILL FILL_1__16963_ (
);

FILL FILL_0__15536_ (
);

AND2X2 _15821_ (
    .A(_4230__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_4770_)
);

FILL FILL_0__15116_ (
);

AND2X2 _15401_ (
    .A(_4189__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_4357_)
);

FILL FILL349600x83980 (
);

FILL FILL94240x133380 (
);

FILL FILL_0__10671_ (
);

FILL FILL472720x103740 (
);

FILL FILL145920x49400 (
);

OR2X2 _18293_ (
    .A(_7204_),
    .B(_7201_),
    .Y(_7205_)
);

FILL FILL131480x335920 (
);

AND2X2 _16606_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_5543_)
);

FILL FILL_0__11876_ (
);

AND2X2 _11741_ (
    .A(_1692_),
    .B(_1691_),
    .Y(_1653_[19])
);

FILL FILL_0__9050_ (
);

FILL FILL66120x266760 (
);

FILL FILL212800x88920 (
);

AND2X2 _11321_ (
    .A(_1472_),
    .B(_1471_),
    .Y(_1455_[8])
);

FILL FILL_0__11036_ (
);

AND2X2 _19498_ (
    .A(_8367_),
    .B(_8366_),
    .Y(_8320_[23])
);

AND2X2 _19078_ (
    .A(_6264__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_7978_)
);

DFFSR _8948_ (
    .CLK(clk_bF$buf85),
    .D(_201_[8]),
    .Q(\datapath_1.regfile_1.regOut[4] [8]),
    .R(rst_bF$buf103),
    .S(vdd)
);

AND2X2 _8528_ (
    .A(_50_),
    .B(_49_),
    .Y(_3_[23])
);

FILL FILL380760x83980 (
);

FILL FILL306280x9880 (
);

FILL FILL441560x24700 (
);

FILL FILL84360x79040 (
);

AND2X2 _12946_ (
    .A(_2509_),
    .B(_2507_),
    .Y(_2510_)
);

FILL FILL_1_BUFX2_insert762 (
);

AND2X2 _12526_ (
    .A(_2115_),
    .B(_2108_),
    .Y(_2116_)
);

OR2X2 _12106_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .B(_1916__bF$buf3),
    .Y(_1876_)
);

FILL FILL_1_BUFX2_insert764 (
);

FILL FILL_1_BUFX2_insert766 (
);

FILL FILL_0__16494_ (
);

FILL FILL_0__16074_ (
);

FILL FILL_1__9631_ (
);

FILL FILL24320x128440 (
);

FILL FILL_1__15814_ (
);

FILL FILL60800x301340 (
);

FILL FILL468920x24700 (
);

FILL FILL_0__14807_ (
);

FILL FILL_1__18286_ (
);

BUFX2 BUFX2_insert430 (
    .A(_6221_),
    .Y(_6221__bF$buf0)
);

BUFX2 BUFX2_insert431 (
    .A(_6315_),
    .Y(_6315__bF$buf4)
);

BUFX2 BUFX2_insert432 (
    .A(_6315_),
    .Y(_6315__bF$buf3)
);

FILL FILL41800x138320 (
);

BUFX2 BUFX2_insert433 (
    .A(_6315_),
    .Y(_6315__bF$buf2)
);

FILL FILL364800x212420 (
);

AND2X2 _17984_ (
    .A(_6321__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_6901_)
);

BUFX2 BUFX2_insert434 (
    .A(_6315_),
    .Y(_6315__bF$buf1)
);

AND2X2 _17564_ (
    .A(_6321__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_6487_)
);

BUFX2 BUFX2_insert435 (
    .A(_6315_),
    .Y(_6315__bF$buf0)
);

BUFX2 BUFX2_insert436 (
    .A(_1124_),
    .Y(_1124__bF$buf4)
);

OR2X2 _17144_ (
    .A(_6072_),
    .B(_6057_),
    .Y(_6073_)
);

BUFX2 BUFX2_insert437 (
    .A(_1124_),
    .Y(_1124__bF$buf3)
);

BUFX2 BUFX2_insert438 (
    .A(_1124_),
    .Y(_1124__bF$buf2)
);

BUFX2 BUFX2_insert439 (
    .A(_1124_),
    .Y(_1124__bF$buf1)
);

FILL FILL_0__18640_ (
);

FILL FILL_0__18220_ (
);

FILL FILL241680x247000 (
);

DFFSR _9486_ (
    .CLK(clk_bF$buf30),
    .D(_465_[30]),
    .Q(\datapath_1.regfile_1.regOut[8] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL451440x123500 (
);

OR2X2 _9066_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_329_)
);

FILL FILL41040x365560 (
);

FILL FILL_0__8741_ (
);

FILL FILL_0__10727_ (
);

FILL FILL_0__10307_ (
);

OR2X2 _18769_ (
    .A(_7673_),
    .B(_7672_),
    .Y(_7674_)
);

FILL FILL90440x163020 (
);

OR2X2 _18349_ (
    .A(_7252_),
    .B(_7259_),
    .Y(_7260_)
);

FILL FILL327560x4940 (
);

FILL FILL250800x0 (
);

FILL FILL_0__13199_ (
);

AND2X2 _13484_ (
    .A(_3012_),
    .B(_3011_),
    .Y(\datapath_1.a3 [3])
);

OR2X2 _13064_ (
    .A(_2387__bF$buf1),
    .B(_2620_),
    .Y(_2621_)
);

FILL FILL_0__19425_ (
);

FILL FILL_0__19005_ (
);

FILL FILL_0__14980_ (
);

FILL FILL_0__14140_ (
);

FILL FILL275880x74100 (
);

FILL FILL_1__12519_ (
);

FILL FILL_0__9946_ (
);

AND2X2 _14689_ (
    .A(_3845_),
    .B(_3844_),
    .Y(_3804_[20])
);

FILL FILL193040x187720 (
);

AND2X2 _14269_ (
    .A(_3625_),
    .B(_3624_),
    .Y(_3606_[9])
);

FILL FILL_0__15765_ (
);

FILL FILL_0__15345_ (
);

AND2X2 _15630_ (
    .A(_4146__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_4582_)
);

AND2X2 _15210_ (
    .A(_4167__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_4168_)
);

FILL FILL_0__10480_ (
);

FILL FILL_0__10060_ (
);

FILL FILL408120x316160 (
);

FILL FILL449920x98800 (
);

OR2X2 _10189_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .B(_926__bF$buf2),
    .Y(_898_)
);

FILL FILL_1__17137_ (
);

FILL FILL_1__12272_ (
);

FILL FILL320720x148200 (
);

AND2X2 _16835_ (
    .A(_4154__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_5768_)
);

OR2X2 _16415_ (
    .A(_5353_),
    .B(_5354_),
    .Y(_5355_)
);

OR2X2 _11970_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_1805_)
);

DFFSR _11550_ (
    .CLK(clk_bF$buf32),
    .D(_1521_[30]),
    .Q(\datapath_1.regfile_1.regOut[24] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

OR2X2 _11130_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_1385_)
);

FILL FILL_0__17911_ (
);

FILL FILL408880x301340 (
);

FILL FILL337440x291460 (
);

FILL FILL256120x227240 (
);

OR2X2 _8757_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_163_)
);

FILL FILL342000x24700 (
);

FILL FILL_1__13477_ (
);

INVX1 _12755_ (
    .A(_2319_),
    .Y(_2320_)
);

AND2X2 _12335_ (
    .A(_1988_),
    .B(_1987_),
    .Y(_1983_[2])
);

FILL FILL_0__13411_ (
);

FILL FILL296400x321100 (
);

FILL FILL87400x316160 (
);

FILL FILL_1__9440_ (
);

FILL FILL37240x167960 (
);

FILL FILL73720x340860 (
);

OR2X2 _14901_ (
    .A(\datapath_1.mux_pcsrc.dout [5]),
    .B(_4001__bF$buf3),
    .Y(_3947_)
);

FILL FILL386080x182780 (
);

FILL FILL9880x301340 (
);

AND2X2 _17793_ (
    .A(_6315__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_6713_)
);

OR2X2 _17373_ (
    .A(_6294_),
    .B(_6298_),
    .Y(_6299_)
);

FILL FILL_0__17088_ (
);

OR2X2 _9295_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .B(_464__bF$buf1),
    .Y(_442_)
);

FILL FILL_1__11963_ (
);

FILL FILL60040x345800 (
);

FILL FILL495520x148200 (
);

FILL FILL_0__8550_ (
);

OR2X2 _10821_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_1219_)
);

FILL FILL_0__10536_ (
);

OR2X2 _10401_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_999_)
);

OR2X2 _18998_ (
    .A(_7891_),
    .B(_7898_),
    .Y(_7899_)
);

OR2X2 _18578_ (
    .A(_7454_),
    .B(_7485_),
    .Y(_7486_)
);

OR2X2 _18158_ (
    .A(_7070_),
    .B(_7071_),
    .Y(_7072_)
);

FILL FILL481840x172900 (
);

FILL FILL383800x74100 (
);

FILL FILL130720x59280 (
);

INVX1 _13293_ (
    .A(_2835_),
    .Y(\datapath_1.ALUResult [9])
);

FILL FILL329840x9880 (
);

FILL FILL_0__19234_ (
);

FILL FILL360240x74100 (
);

FILL FILL134520x360620 (
);

FILL FILL_1__12328_ (
);

FILL FILL504640x118560 (
);

FILL FILL_0__9755_ (
);

AND2X2 _11606_ (
    .A(_1622_),
    .B(_1621_),
    .Y(_1587_[17])
);

FILL FILL320720x375440 (
);

INVX2 _14498_ (
    .A(IRWrite_bF$buf4),
    .Y(_3803_)
);

OR2X2 _14078_ (
    .A(_3486_),
    .B(_3483_),
    .Y(\datapath_1.alu_1.ALUInB [22])
);

FILL FILL_0__15994_ (
);

FILL FILL_0__15574_ (
);

FILL FILL161880x316160 (
);

FILL FILL_1__17786_ (
);

FILL FILL367840x9880 (
);

FILL FILL_1__17366_ (
);

FILL FILL269800x360620 (
);

OR2X2 _16644_ (
    .A(_5579_),
    .B(_5578_),
    .Y(_5580_)
);

FILL FILL_0__16359_ (
);

OR2X2 _16224_ (
    .A(_5163_),
    .B(_5166_),
    .Y(_5167_)
);

FILL FILL_0__11494_ (
);

FILL FILL_0__17300_ (
);

OR2X2 _8986_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_332__bF$buf4),
    .Y(_276_)
);

DFFSR _8566_ (
    .CLK(clk_bF$buf47),
    .D(_3_[13]),
    .Q(\datapath_1.regfile_1.regOut[1] [13]),
    .R(rst_bF$buf103),
    .S(vdd)
);

OR2X2 _17849_ (
    .A(_6766_),
    .B(_6767_),
    .Y(_6768_)
);

FILL FILL286520x276640 (
);

NOR2X1 _17429_ (
    .A(_6310__bF$buf3),
    .B(_6353_),
    .Y(_6354_)
);

AND2X2 _17009_ (
    .A(_4183__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_5940_)
);

FILL FILL_0__12699_ (
);

XOR2X1 _12984_ (
    .A(_2325_),
    .B(_2544_),
    .Y(_2545_)
);

NOR2X1 _12564_ (
    .A(_2111_),
    .B(_2133_),
    .Y(_2085_)
);

OR2X2 _12144_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_1901_)
);

FILL FILL381520x98800 (
);

FILL FILL392160x350740 (
);

FILL FILL_0__18925_ (
);

FILL FILL_0__18505_ (
);

FILL FILL_0__13640_ (
);

FILL FILL132240x222300 (
);

FILL FILL_0__8606_ (
);

AND2X2 _13769_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [25]),
    .Y(_3239_)
);

AND2X2 _13349_ (
    .A(_2888_),
    .B(_2880_),
    .Y(_2889_)
);

FILL FILL_1__15432_ (
);

AND2X2 _14710_ (
    .A(_3859_),
    .B(_3858_),
    .Y(_3804_[27])
);

FILL FILL_0__14425_ (
);

FILL FILL_0__14005_ (
);

BUFX2 BUFX2_insert810 (
    .A(_6323_),
    .Y(_6323__bF$buf2)
);

BUFX2 BUFX2_insert811 (
    .A(_6323_),
    .Y(_6323__bF$buf1)
);

BUFX2 BUFX2_insert812 (
    .A(_6323_),
    .Y(_6323__bF$buf0)
);

BUFX2 BUFX2_insert813 (
    .A(_6264_),
    .Y(_6264__bF$buf4)
);

BUFX2 BUFX2_insert814 (
    .A(_6264_),
    .Y(_6264__bF$buf3)
);

BUFX2 BUFX2_insert815 (
    .A(_6264_),
    .Y(_6264__bF$buf2)
);

BUFX2 BUFX2_insert816 (
    .A(_6264_),
    .Y(_6264__bF$buf1)
);

AND2X2 _17182_ (
    .A(_4142__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_6110_)
);

BUFX2 BUFX2_insert817 (
    .A(_6264_),
    .Y(_6264__bF$buf0)
);

BUFX2 BUFX2_insert818 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf4 )
);

BUFX2 BUFX2_insert819 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf3 )
);

FILL FILL350360x212420 (
);

FILL FILL385320x98800 (
);

FILL FILL_1__11772_ (
);

OR2X2 _15915_ (
    .A(_4862_),
    .B(_4861_),
    .Y(_4863_)
);

FILL FILL267520x222300 (
);

DFFSR _10630_ (
    .CLK(clk_bF$buf63),
    .D(_1059_[13]),
    .Q(\datapath_1.regfile_1.regOut[17] [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

OR2X2 _10210_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_926__bF$buf2),
    .Y(_912_)
);

AND2X2 _18387_ (
    .A(_6312__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_7297_)
);

FILL FILL278920x291460 (
);

FILL FILL468160x202540 (
);

FILL FILL_0__9564_ (
);

OR2X2 _11835_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_1735_)
);

FILL FILL_0__9144_ (
);

DFFSR _11415_ (
    .CLK(clk_bF$buf96),
    .D(_1455_[24]),
    .Q(\datapath_1.regfile_1.regOut[23] [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL_0__12911_ (
);

FILL FILL398240x207480 (
);

FILL FILL_1__16390_ (
);

FILL FILL265240x296400 (
);

FILL FILL_0__15383_ (
);

FILL FILL475000x172900 (
);

FILL FILL_1__8520_ (
);

FILL FILL208240x64220 (
);

FILL FILL_0__16588_ (
);

AND2X2 _16873_ (
    .A(_4203__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_5806_)
);

AND2X2 _16453_ (
    .A(_4217__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_5392_)
);

AND2X2 _16033_ (
    .A(_4230__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_4979_)
);

AND2X2 _8795_ (
    .A(_188_),
    .B(_187_),
    .Y(_135_[26])
);

FILL FILL_1__15908_ (
);

FILL FILL272840x232180 (
);

FILL FILL141360x340860 (
);

FILL FILL_1__13095_ (
);

OR2X2 _17658_ (
    .A(_6579_),
    .B(_6576_),
    .Y(_6580_)
);

OR2X2 _17238_ (
    .A(_6163_),
    .B(_6164_),
    .Y(_6165_)
);

OR2X2 _12793_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2358_)
);

OR2X2 _12373_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .B(_2048__bF$buf1),
    .Y(_2014_)
);

FILL FILL436240x14820 (
);

FILL FILL_0__18734_ (
);

FILL FILL259920x103740 (
);

FILL FILL_0__8415_ (
);

FILL FILL6840x158080 (
);

AND2X2 _13998_ (
    .A(_3350__bF$buf2),
    .B(_2_[11]),
    .Y(_3418_)
);

AND2X2 _13578_ (
    .A(_3073_),
    .B(_3072_),
    .Y(_1_[29])
);

NAND2X1 _13158_ (
    .A(_2696_),
    .B(_2708_),
    .Y(_2709_)
);

FILL FILL139080x49400 (
);

FILL FILL_0__19519_ (
);

FILL FILL_0__14654_ (
);

FILL FILL_0__14234_ (
);

FILL FILL380000x276640 (
);

FILL FILL413440x88920 (
);

FILL FILL449920x360620 (
);

FILL FILL_1__11581_ (
);

FILL FILL_0__15859_ (
);

FILL FILL_0__15439_ (
);

AND2X2 _15724_ (
    .A(_4228__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_4675_)
);

OR2X2 _15304_ (
    .A(_4257_),
    .B(_4260_),
    .Y(_4261_)
);

FILL FILL202920x227240 (
);

FILL FILL_0__10994_ (
);

FILL FILL_0__10574_ (
);

FILL FILL293360x256880 (
);

OR2X2 _18196_ (
    .A(_7108_),
    .B(_7107_),
    .Y(_7109_)
);

FILL FILL63080x261820 (
);

FILL FILL_0__16800_ (
);

FILL FILL_0__19272_ (
);

AND2X2 _16929_ (
    .A(_4151__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_5861_)
);

OR2X2 _16509_ (
    .A(_5445_),
    .B(_5446_),
    .Y(_5447_)
);

FILL FILL_0__9373_ (
);

OR2X2 _11644_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .B(_1652__bF$buf4),
    .Y(_1648_)
);

OR2X2 _11224_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .B(_1454__bF$buf4),
    .Y(_1428_)
);

FILL FILL53960x74100 (
);

FILL FILL_0__15192_ (
);

AND2X2 _12849_ (
    .A(_2409_),
    .B(_2413_),
    .Y(_2414_)
);

DFFSR _12429_ (
    .CLK(clk_bF$buf49),
    .D(_1983_[6]),
    .Q(\datapath_1.regfile_1.regOut[31] [6]),
    .R(rst_bF$buf106),
    .S(vdd)
);

OR2X2 _12009_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_1831_)
);

FILL FILL_0__13925_ (
);

FILL FILL_0__13505_ (
);

AND2X2 _16682_ (
    .A(_4142__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_5618_)
);

AND2X2 _16262_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_5204_)
);

FILL FILL_1__9534_ (
);

FILL FILL255360x360620 (
);

FILL FILL74480x24700 (
);

FILL FILL_1__10852_ (
);

FILL FILL82840x207480 (
);

FILL FILL185440x365560 (
);

AND2X2 _17887_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_6805_)
);

AND2X2 _17467_ (
    .A(_6236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_6392_)
);

OR2X2 _17047_ (
    .A(_5976_),
    .B(_5973_),
    .Y(_5977_)
);

DFFSR _12182_ (
    .CLK(clk_bF$buf65),
    .D(_1851_[17]),
    .Q(\datapath_1.regfile_1.regOut[29] [17]),
    .R(rst_bF$buf36),
    .S(vdd)
);

FILL FILL_0__18123_ (
);

AND2X2 _9389_ (
    .A(_484_),
    .B(_483_),
    .Y(_465_[9])
);

FILL FILL272080x276640 (
);

FILL FILL_1__11217_ (
);

FILL FILL_0__8644_ (
);

OR2X2 _10915_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .B(_1322__bF$buf1),
    .Y(_1262_)
);

FILL FILL189240x286520 (
);

NAND3X1 _13387_ (
    .A(_2379__bF$buf2),
    .B(\datapath_1.alu_1.ALUInB [3]),
    .C(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2924_)
);

FILL FILL268280x88920 (
);

FILL FILL263720x24700 (
);

FILL FILL_0__9009_ (
);

FILL FILL405080x311220 (
);

FILL FILL133000x187720 (
);

FILL FILL_1__16255_ (
);

AND2X2 _15953_ (
    .A(_4189__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_4900_)
);

AND2X2 _15533_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_4487_)
);

AND2X2 _15113_ (
    .A(_4092_),
    .B(_4036_),
    .Y(_4093_)
);

FILL FILL166440x311220 (
);

FILL FILL_1__8805_ (
);

FILL FILL253080x222300 (
);

FILL FILL3800x192660 (
);

FILL FILL_1__12595_ (
);

AND2X2 _16738_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_5673_)
);

AND2X2 _16318_ (
    .A(_4151__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_5259_)
);

FILL FILL_0__11588_ (
);

AND2X2 _11873_ (
    .A(_1760_),
    .B(_1759_),
    .Y(_1719_[20])
);

FILL FILL_0__9182_ (
);

AND2X2 _11453_ (
    .A(_1540_),
    .B(_1539_),
    .Y(_1521_[9])
);

FILL FILL_0__11168_ (
);

DFFSR _11033_ (
    .CLK(clk_bF$buf53),
    .D(_1257_[29]),
    .Q(\datapath_1.regfile_1.regOut[20] [29]),
    .R(rst_bF$buf31),
    .S(vdd)
);

FILL FILL_0__17814_ (
);

FILL FILL_1__10908_ (
);

DFFSR _9601_ (
    .CLK(clk_bF$buf5),
    .D(_531_[16]),
    .Q(\datapath_1.regfile_1.regOut[9] [16]),
    .R(rst_bF$buf10),
    .S(vdd)
);

NAND2X1 _12658_ (
    .A(_2221_),
    .B(_2222_),
    .Y(_2223_)
);

OR2X2 _12238_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .B(_1982__bF$buf2),
    .Y(_1944_)
);

FILL FILL_0__13734_ (
);

FILL FILL_0_BUFX2_insert1150 (
);

FILL FILL_0_BUFX2_insert1151 (
);

FILL FILL_0_BUFX2_insert1152 (
);

OR2X2 _16491_ (
    .A(_5429_),
    .B(_5428_),
    .Y(_5430_)
);

FILL FILL_0_BUFX2_insert1154 (
);

OR2X2 _16071_ (
    .A(_5014_),
    .B(_5015_),
    .Y(_5016_)
);

FILL FILL_0_BUFX2_insert1156 (
);

FILL FILL_0_BUFX2_insert1158 (
);

FILL FILL_1__10661_ (
);

FILL FILL_0__14939_ (
);

OR2X2 _14804_ (
    .A(vdd),
    .B(_2_[16]),
    .Y(_3902_)
);

FILL FILL_0__14519_ (
);

FILL FILL152760x158080 (
);

FILL FILL437000x301340 (
);

AND2X2 _17696_ (
    .A(_6264__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_6617_)
);

INVX1 _17276_ (
    .A(\datapath_1.PCJump [24]),
    .Y(_6202_)
);

FILL FILL_0__18772_ (
);

FILL FILL_0__18352_ (
);

DFFSR _9198_ (
    .CLK(clk_bF$buf41),
    .D(_333_[0]),
    .Q(\datapath_1.regfile_1.regOut[6] [0]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL99560x167960 (
);

FILL FILL_0__8873_ (
);

FILL FILL_0__8453_ (
);

FILL FILL_0__10859_ (
);

FILL FILL_0__10439_ (
);

AND2X2 _10724_ (
    .A(_1174_),
    .B(_1173_),
    .Y(_1125_[24])
);

FILL FILL_0__10019_ (
);

AND2X2 _10304_ (
    .A(_954_),
    .B(_953_),
    .Y(_927_[13])
);

OR2X2 _13196_ (
    .A(_2421_),
    .B(_2744_),
    .Y(_2745_)
);

FILL FILL_0__19557_ (
);

OR2X2 _19422_ (
    .A(_8301_),
    .B(_8316_),
    .Y(_8317_)
);

FILL FILL_0__19137_ (
);

AND2X2 _19002_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_7903_)
);

FILL FILL175560x108680 (
);

FILL FILL_0__14692_ (
);

FILL FILL57760x163020 (
);

FILL FILL_0__9658_ (
);

DFFSR _11929_ (
    .CLK(clk_bF$buf101),
    .D(_1719_[22]),
    .Q(\datapath_1.regfile_1.regOut[27] [22]),
    .R(rst_bF$buf54),
    .S(vdd)
);

OR2X2 _11509_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .B(_1586__bF$buf3),
    .Y(_1578_)
);

FILL FILL_1__16484_ (
);

AND2X2 _15762_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_4712_)
);

FILL FILL_0__15477_ (
);

FILL FILL_0__15057_ (
);

OR2X2 _15342_ (
    .A(_4297_),
    .B(_4298_),
    .Y(_4299_)
);

FILL FILL_0__10192_ (
);

FILL FILL29640x296400 (
);

FILL FILL416480x197600 (
);

FILL FILL260680x187720 (
);

OR2X2 _16967_ (
    .A(_5897_),
    .B(_5896_),
    .Y(_5898_)
);

OR2X2 _16547_ (
    .A(_5484_),
    .B(_5483_),
    .Y(_5485_)
);

AND2X2 _16127_ (
    .A(_4172__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_5071_)
);

INVX2 _11682_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .Y(_1718_)
);

DFFSR _11262_ (
    .CLK(clk_bF$buf19),
    .D(_1389_[0]),
    .Q(\datapath_1.regfile_1.regOut[22] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL_0__17623_ (
);

FILL FILL_0__17203_ (
);

FILL FILL397480x340860 (
);

OR2X2 _8889_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_231_)
);

OR2X2 _8469_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_11_)
);

AND2X2 _9830_ (
    .A(_718_),
    .B(_717_),
    .Y(_663_[27])
);

AND2X2 _9410_ (
    .A(_498_),
    .B(_497_),
    .Y(_465_[16])
);

OR2X2 _12887_ (
    .A(_2450_),
    .B(_2451_),
    .Y(_2452_)
);

FILL FILL_1__19415_ (
);

INVX1 _12467_ (
    .A(\aluControl_1.inst [0]),
    .Y(_2060_)
);

DFFSR _12047_ (
    .CLK(clk_bF$buf51),
    .D(_1785_[11]),
    .Q(\datapath_1.regfile_1.regOut[28] [11]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL_1__14970_ (
);

FILL FILL_0__13963_ (
);

FILL FILL_0__13543_ (
);

FILL FILL_0__13123_ (
);

FILL FILL505400x370500 (
);

FILL FILL_0__8929_ (
);

FILL FILL_1__9572_ (
);

FILL FILL122360x79040 (
);

FILL FILL_0__14328_ (
);

DFFSR _14613_ (
    .CLK(clk_bF$buf65),
    .D(_3738_[19]),
    .Q(\datapath_1.PCJump [21]),
    .R(rst_bF$buf26),
    .S(vdd)
);

FILL FILL171760x138320 (
);

OR2X2 _17085_ (
    .A(_6013_),
    .B(_6012_),
    .Y(_6014_)
);

FILL FILL129960x64220 (
);

AND2X2 _15818_ (
    .A(_4175__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_4767_)
);

FILL FILL493240x291460 (
);

FILL FILL149720x79040 (
);

OR2X2 _10953_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_1287_)
);

FILL FILL_0__10668_ (
);

OR2X2 _10533_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_1067_)
);

DFFSR _10113_ (
    .CLK(clk_bF$buf102),
    .D(_795_[12]),
    .Q(\datapath_1.regfile_1.regOut[13] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

FILL FILL292600x177840 (
);

FILL FILL102600x49400 (
);

FILL FILL_0__19366_ (
);

AND2X2 _19231_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_8128_)
);

FILL FILL_0__14081_ (
);

FILL FILL132240x182780 (
);

FILL FILL_0__9887_ (
);

FILL FILL123880x88920 (
);

AND2X2 _11738_ (
    .A(_1690_),
    .B(_1689_),
    .Y(_1653_[18])
);

FILL FILL_0__9047_ (
);

AND2X2 _11318_ (
    .A(_1470_),
    .B(_1469_),
    .Y(_1455_[7])
);

FILL FILL357960x14820 (
);

FILL FILL_1__13401_ (
);

OR2X2 _15991_ (
    .A(_4930_),
    .B(_4937_),
    .Y(_4938_)
);

OR2X2 _15571_ (
    .A(_4523_),
    .B(_4522_),
    .Y(_4524_)
);

OAI21X1 _15151_ (
    .A(_4005_),
    .B(_4094_),
    .C(\datapath_1.a3 [4]),
    .Y(_4116_)
);

FILL FILL21280x64220 (
);

FILL FILL38000x217360 (
);

OR2X2 _16776_ (
    .A(_5706_),
    .B(_5709_),
    .Y(_5710_)
);

AND2X2 _16356_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_5297_)
);

FILL FILL273600x123500 (
);

OR2X2 _11491_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .B(_1586__bF$buf3),
    .Y(_1566_)
);

OR2X2 _11071_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .B(_1388__bF$buf2),
    .Y(_1346_)
);

FILL FILL_0__17852_ (
);

FILL FILL_0__17012_ (
);

FILL FILL465120x212420 (
);

DFFSR _8698_ (
    .CLK(clk_bF$buf64),
    .D(_69_[16]),
    .Q(\datapath_1.regfile_1.regOut[2] [16]),
    .R(rst_bF$buf10),
    .S(vdd)
);

FILL FILL212800x232180 (
);

FILL FILL19760x360620 (
);

FILL FILL210520x64220 (
);

FILL FILL32680x355680 (
);

INVX1 _12696_ (
    .A(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2261_)
);

OR2X2 _12276_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_1969_)
);

FILL FILL_0__18637_ (
);

AND2X2 _18922_ (
    .A(_6247__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_7824_)
);

FILL FILL_0__18217_ (
);

OR2X2 _18502_ (
    .A(_7410_),
    .B(_7409_),
    .Y(_7411_)
);

FILL FILL_0__13352_ (
);

FILL FILL271320x197600 (
);

FILL FILL_0__8738_ (
);

FILL FILL359480x350740 (
);

FILL FILL_1__9381_ (
);

FILL FILL_1__15984_ (
);

FILL FILL_0__14977_ (
);

AND2X2 _14842_ (
    .A(_3927_),
    .B(_3926_),
    .Y(_3870_[28])
);

FILL FILL_0__14557_ (
);

AND2X2 _14422_ (
    .A(_3707_),
    .B(_3706_),
    .Y(_3672_[17])
);

AND2X2 _14002_ (
    .A(_3344__bF$buf0),
    .B(gnd),
    .Y(_3421_)
);

FILL FILL395960x79040 (
);

FILL FILL69160x14820 (
);

FILL FILL429400x24700 (
);

FILL FILL30400x326040 (
);

FILL FILL164920x49400 (
);

FILL FILL_0__18390_ (
);

FILL FILL_1__16769_ (
);

FILL FILL_1__16349_ (
);

FILL FILL345040x83980 (
);

AND2X2 _15627_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_4579_)
);

AND2X2 _15207_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_4165_)
);

FILL FILL13680x301340 (
);

FILL FILL_0__8491_ (
);

DFFSR _10762_ (
    .CLK(clk_bF$buf76),
    .D(_1125_[16]),
    .Q(\datapath_1.regfile_1.regOut[18] [16]),
    .R(rst_bF$buf112),
    .S(vdd)
);

OR2X2 _10342_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .B(_992__bF$buf3),
    .Y(_980_)
);

AND2X2 _18099_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_7014_)
);

FILL FILL389880x172900 (
);

FILL FILL317680x212420 (
);

FILL FILL_0__19175_ (
);

OR2X2 _19460_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_8342_)
);

AND2X2 _19040_ (
    .A(_6293__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [26]),
    .Y(_7940_)
);

FILL FILL20520x271700 (
);

OR2X2 _8910_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_245_)
);

FILL FILL_0__9696_ (
);

OR2X2 _11967_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_1803_)
);

FILL FILL_0__9276_ (
);

DFFSR _11547_ (
    .CLK(clk_bF$buf68),
    .D(_1521_[27]),
    .Q(\datapath_1.regfile_1.regOut[24] [27]),
    .R(rst_bF$buf40),
    .S(vdd)
);

OR2X2 _11127_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_1383_)
);

FILL FILL_0__12623_ (
);

FILL FILL_0__12203_ (
);

FILL FILL236360x74100 (
);

FILL FILL168720x49400 (
);

FILL FILL_0__15095_ (
);

AND2X2 _15380_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_4336_)
);

FILL FILL133760x335920 (
);

FILL FILL_1__8652_ (
);

FILL FILL_1__14415_ (
);

FILL FILL465880x207480 (
);

FILL FILL_0__13828_ (
);

FILL FILL_0__13408_ (
);

FILL FILL455240x167960 (
);

OR2X2 _16585_ (
    .A(_5514_),
    .B(_5521_),
    .Y(_5522_)
);

AND2X2 _16165_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_5109_)
);

FILL FILL491720x340860 (
);

FILL FILL_0__17241_ (
);

FILL FILL_1__19033_ (
);

OR2X2 _12085_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_1916__bF$buf2),
    .Y(_1862_)
);

FILL FILL_0__18866_ (
);

FILL FILL222680x316160 (
);

OR2X2 _18731_ (
    .A(_7632_),
    .B(_7635_),
    .Y(_7636_)
);

FILL FILL_0__18446_ (
);

OR2X2 _18311_ (
    .A(_7221_),
    .B(_7222_),
    .Y(_7223_)
);

FILL FILL_0__13581_ (
);

FILL FILL212040x276640 (
);

FILL FILL139840x326040 (
);

FILL FILL26600x128440 (
);

FILL FILL_0__8547_ (
);

OR2X2 _10818_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_1217_)
);

FILL FILL_1__12901_ (
);

FILL FILL_1__15373_ (
);

AND2X2 _19516_ (
    .A(_8379_),
    .B(_8378_),
    .Y(_8320_[29])
);

FILL FILL_0__14786_ (
);

OR2X2 _14651_ (
    .A(vdd),
    .B(\datapath_1.a [8]),
    .Y(_3820_)
);

OR2X2 _14231_ (
    .A(\datapath_1.Data [29]),
    .B(_3605__bF$buf0),
    .Y(_3599_)
);

FILL FILL468160x24700 (
);

FILL FILL252320x370500 (
);

FILL FILL453720x123500 (
);

FILL FILL_1__16998_ (
);

FILL FILL92720x163020 (
);

AND2X2 _15856_ (
    .A(_4236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_4805_)
);

OR2X2 _15436_ (
    .A(_4389_),
    .B(_4390_),
    .Y(_4391_)
);

INVX1 _15016_ (
    .A(\datapath_1.a3 [3]),
    .Y(_4005_)
);

AND2X2 _10991_ (
    .A(_1312_),
    .B(_1311_),
    .Y(_1257_[27])
);

AND2X2 _10571_ (
    .A(_1092_),
    .B(_1091_),
    .Y(_1059_[16])
);

AND2X2 _10151_ (
    .A(_872_),
    .B(_871_),
    .Y(_861_[5])
);

FILL FILL_0__16932_ (
);

FILL FILL_0__16512_ (
);

FILL FILL445360x98800 (
);

FILL FILL_1__12078_ (
);

OR2X2 _11776_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .B(_1718__bF$buf0),
    .Y(_1716_)
);

OR2X2 _11356_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .B(_1520__bF$buf4),
    .Y(_1496_)
);

FILL FILL_0__17717_ (
);

FILL FILL_0__12852_ (
);

FILL FILL_0__12012_ (
);

OR2X2 _9924_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_761_)
);

OR2X2 _9504_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_541_)
);

FILL FILL_1__8461_ (
);

FILL FILL_1__19509_ (
);

FILL FILL_1__14224_ (
);

FILL FILL240920x330980 (
);

FILL FILL328320x222300 (
);

AND2X2 _13922_ (
    .A(_3352__bF$buf4),
    .B(gnd),
    .Y(_3353_)
);

FILL FILL_0__13217_ (
);

OR2X2 _13502_ (
    .A(ALUOut[4]),
    .B(_3079__bF$buf3),
    .Y(_3023_)
);

FILL FILL422560x281580 (
);

FILL FILL47880x29640 (
);

FILL FILL104880x370500 (
);

AND2X2 _16394_ (
    .A(_4203__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_5334_)
);

FILL FILL339720x291460 (
);

FILL FILL_1__9666_ (
);

FILL FILL_0__17890_ (
);

FILL FILL_0__17470_ (
);

FILL FILL_1__15849_ (
);

FILL FILL_1__10984_ (
);

AND2X2 _14707_ (
    .A(_3857_),
    .B(_3856_),
    .Y(_3804_[26])
);

BUFX2 BUFX2_insert780 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf2 )
);

BUFX2 BUFX2_insert781 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf1 )
);

BUFX2 BUFX2_insert782 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf0 )
);

BUFX2 BUFX2_insert783 (
    .A(_4142_),
    .Y(_4142__bF$buf4)
);

BUFX2 BUFX2_insert784 (
    .A(_4142_),
    .Y(_4142__bF$buf3)
);

OR2X2 _17599_ (
    .A(_6520_),
    .B(_6521_),
    .Y(_6522_)
);

BUFX2 BUFX2_insert785 (
    .A(_4142_),
    .Y(_4142__bF$buf2)
);

BUFX2 BUFX2_insert786 (
    .A(_4142_),
    .Y(_4142__bF$buf1)
);

AND2X2 _17179_ (
    .A(_4130__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_6107_)
);

BUFX2 BUFX2_insert787 (
    .A(_4142_),
    .Y(_4142__bF$buf0)
);

BUFX2 BUFX2_insert788 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf4 )
);

BUFX2 BUFX2_insert789 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf3 )
);

AND2X2 _18960_ (
    .A(_6300__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_7862_)
);

FILL FILL_0__18255_ (
);

AND2X2 _18540_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_7448_)
);

OR2X2 _18120_ (
    .A(_7031_),
    .B(_7034_),
    .Y(_7035_)
);

FILL FILL408880x375440 (
);

FILL FILL_1__11349_ (
);

FILL FILL_0__8776_ (
);

DFFSR _10627_ (
    .CLK(clk_bF$buf30),
    .D(_1059_[10]),
    .Q(\datapath_1.regfile_1.regOut[17] [10]),
    .R(rst_bF$buf84),
    .S(vdd)
);

OR2X2 _10207_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .B(_926__bF$buf0),
    .Y(_910_)
);

INVX1 _13099_ (
    .A(_2653_),
    .Y(\datapath_1.ALUResult [21])
);

FILL FILL_0__11703_ (
);

OR2X2 _19325_ (
    .A(_8220_),
    .B(_8207_),
    .Y(_8221_)
);

FILL FILL117040x69160 (
);

DFFSR _14880_ (
    .CLK(clk_bF$buf98),
    .D(_3870_[28]),
    .Q(_2_[28]),
    .R(rst_bF$buf87),
    .S(vdd)
);

FILL FILL_0__14175_ (
);

OR2X2 _14460_ (
    .A(memoryOutData[30]),
    .B(_3737__bF$buf0),
    .Y(_3733_)
);

AND2X2 _14040_ (
    .A(_3350__bF$buf0),
    .B(_2_[17]),
    .Y(_3454_)
);

FILL FILL10640x158080 (
);

FILL FILL333640x232180 (
);

FILL FILL202160x340860 (
);

FILL FILL_0__12908_ (
);

FILL FILL420280x143260 (
);

AND2X2 _15665_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_4617_)
);

AND2X2 _15245_ (
    .A(_4202_),
    .B(_4144_),
    .Y(_4203_)
);

DFFSR _10380_ (
    .CLK(clk_bF$buf21),
    .D(_927_[21]),
    .Q(\datapath_1.regfile_1.regOut[15] [21]),
    .R(rst_bF$buf90),
    .S(vdd)
);

FILL FILL_1__8937_ (
);

FILL FILL_0__16741_ (
);

FILL FILL_0__16321_ (
);

FILL FILL136800x360620 (
);

FILL FILL181640x143260 (
);

FILL FILL_1__18533_ (
);

AND2X2 _11585_ (
    .A(_1608_),
    .B(_1607_),
    .Y(_1587_[10])
);

FILL FILL_1__18113_ (
);

OR2X2 _11165_ (
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .Y(_1453_)
);

OR2X2 _17811_ (
    .A(_6729_),
    .B(_6728_),
    .Y(_6730_)
);

FILL FILL_0__17106_ (
);

FILL FILL_0__12661_ (
);

FILL FILL_0__12241_ (
);

DFFSR _9733_ (
    .CLK(clk_bF$buf60),
    .D(_597_[19]),
    .Q(\datapath_1.regfile_1.regOut[10] [19]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9313_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .B(_464__bF$buf2),
    .Y(_454_)
);

FILL FILL424080x251940 (
);

FILL FILL28880x227240 (
);

FILL FILL_0__13446_ (
);

AND2X2 _13731_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[20]),
    .Y(_3206_)
);

XNOR2X1 _13311_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2852_)
);

FILL FILL_1__15238_ (
);

FILL FILL_1__10793_ (
);

FILL FILL199880x212420 (
);

OR2X2 _14936_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [17]),
    .Y(_3970_)
);

OR2X2 _14516_ (
    .A(IRWrite_bF$buf3),
    .B(\datapath_1.PCJump [8]),
    .Y(_3750_)
);

FILL FILL_0__18484_ (
);

FILL FILL205200x54340 (
);

FILL FILL_0__18064_ (
);

FILL FILL433960x93860 (
);

FILL FILL134520x222300 (
);

FILL FILL504640x301340 (
);

FILL FILL_0__8585_ (
);

AND2X2 _10856_ (
    .A(_1242_),
    .B(_1241_),
    .Y(_1191_[25])
);

AND2X2 _10436_ (
    .A(_1022_),
    .B(_1021_),
    .Y(_993_[14])
);

AND2X2 _10016_ (
    .A(_802_),
    .B(_801_),
    .Y(_795_[3])
);

FILL FILL_0__11512_ (
);

FILL FILL12160x128440 (
);

DFFSR _19554_ (
    .CLK(clk_bF$buf9),
    .D(_8320_[31]),
    .Q(\datapath_1.regfile_1.regOut[0] [31]),
    .R(rst_bF$buf23),
    .S(vdd)
);

AND2X2 _19134_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_8033_)
);

FILL FILL_1__13724_ (
);

FILL FILL_0__12717_ (
);

FILL FILL269800x222300 (
);

FILL FILL46360x281580 (
);

OR2X2 _15894_ (
    .A(_4841_),
    .B(_4840_),
    .Y(_4842_)
);

OR2X2 _15474_ (
    .A(_4427_),
    .B(_4428_),
    .Y(_4429_)
);

FILL FILL_0__15189_ (
);

INVX1 _15054_ (
    .A(_4042_),
    .Y(_4043_)
);

FILL FILL89680x345800 (
);

FILL FILL_0__16970_ (
);

OR2X2 _16679_ (
    .A(_5614_),
    .B(_5611_),
    .Y(_5615_)
);

AND2X2 _16259_ (
    .A(_4236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_5201_)
);

FILL FILL_1__18762_ (
);

DFFSR _11394_ (
    .CLK(clk_bF$buf100),
    .D(_1455_[3]),
    .Q(\datapath_1.regfile_1.regOut[23] [3]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL267520x296400 (
);

FILL FILL_0__17755_ (
);

OR2X2 _17620_ (
    .A(_6541_),
    .B(_6537_),
    .Y(_6542_)
);

FILL FILL_0__17335_ (
);

AND2X2 _17200_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_6128_)
);

FILL FILL_0__12470_ (
);

FILL FILL_1__10009_ (
);

AND2X2 _9962_ (
    .A(_786_),
    .B(_785_),
    .Y(_729_[28])
);

AND2X2 _9542_ (
    .A(_566_),
    .B(_565_),
    .Y(_531_[17])
);

AND2X2 _9122_ (
    .A(_346_),
    .B(_345_),
    .Y(_333_[6])
);

INVX1 _12599_ (
    .A(\datapath_1.alu_1.ALUInA [30]),
    .Y(_2164_)
);

DFFSR _12179_ (
    .CLK(clk_bF$buf22),
    .D(_1851_[14]),
    .Q(\datapath_1.regfile_1.regOut[29] [14]),
    .R(rst_bF$buf7),
    .S(vdd)
);

AND2X2 _18825_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_7729_)
);

FILL FILL_0_BUFX2_insert421 (
);

OR2X2 _18405_ (
    .A(_7311_),
    .B(_7314_),
    .Y(_7315_)
);

FILL FILL_0_BUFX2_insert423 (
);

AND2X2 _13960_ (
    .A(_3344__bF$buf3),
    .B(gnd),
    .Y(_3385_)
);

FILL FILL_0__13675_ (
);

OR2X2 _13540_ (
    .A(IorD_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [17]),
    .Y(_3048_)
);

FILL FILL_0_BUFX2_insert425 (
);

NOR2X1 _13120_ (
    .A(_2278_),
    .B(_2498_),
    .Y(_2673_)
);

FILL FILL_0_BUFX2_insert426 (
);

FILL FILL_0_BUFX2_insert427 (
);

FILL FILL_0_BUFX2_insert428 (
);

FILL FILL_0_BUFX2_insert429 (
);

FILL FILL485640x286520 (
);

FILL FILL157320x316160 (
);

FILL FILL50920x64220 (
);

FILL FILL_1__15467_ (
);

FILL FILL174800x326040 (
);

FILL FILL58520x24700 (
);

DFFSR _14745_ (
    .CLK(clk_bF$buf94),
    .D(_3804_[22]),
    .Q(\datapath_1.a [22]),
    .R(rst_bF$buf61),
    .S(vdd)
);

OR2X2 _14325_ (
    .A(\datapath_1.ALUResult [28]),
    .B(_3671__bF$buf4),
    .Y(_3663_)
);

FILL FILL_0__15401_ (
);

FILL FILL_0__18293_ (
);

FILL FILL471200x113620 (
);

FILL FILL_0__8394_ (
);

FILL FILL_1__17613_ (
);

OR2X2 _10665_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_1135_)
);

DFFSR _10245_ (
    .CLK(clk_bF$buf89),
    .D(_861_[15]),
    .Q(\datapath_1.regfile_1.regOut[14] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL_0__16606_ (
);

FILL FILL_0__11741_ (
);

FILL FILL_0__11321_ (
);

OR2X2 _19363_ (
    .A(_8256_),
    .B(_8257_),
    .Y(_8258_)
);

FILL FILL_0__19078_ (
);

FILL FILL101840x202540 (
);

DFFSR _8813_ (
    .CLK(clk_bF$buf112),
    .D(_135_[2]),
    .Q(\datapath_1.regfile_1.regOut[3] [2]),
    .R(rst_bF$buf3),
    .S(vdd)
);

FILL FILL92720x326040 (
);

FILL FILL12160x98800 (
);

FILL FILL475000x69160 (
);

FILL FILL396720x237120 (
);

FILL FILL_0__12946_ (
);

OR2X2 _12811_ (
    .A(_2375_),
    .B(_2374_),
    .Y(_2376_)
);

FILL FILL265240x345800 (
);

FILL FILL295640x256880 (
);

FILL FILL65360x261820 (
);

AND2X2 _15283_ (
    .A(_4213_),
    .B(\datapath_1.PCJump_22_bF$buf0 ),
    .Y(_4241_)
);

FILL FILL96520x247000 (
);

OR2X2 _16488_ (
    .A(_5419_),
    .B(_5426_),
    .Y(_5427_)
);

OR2X2 _16068_ (
    .A(_5011_),
    .B(_5012_),
    .Y(_5013_)
);

FILL FILL_0__17984_ (
);

FILL FILL_0__17564_ (
);

FILL FILL497040x79040 (
);

OR2X2 _9771_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_679_)
);

DFFSR _9351_ (
    .CLK(clk_bF$buf97),
    .D(_399_[24]),
    .Q(\datapath_1.regfile_1.regOut[7] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL_0__18769_ (
);

AND2X2 _18634_ (
    .A(_6300__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_7541_)
);

AND2X2 _18214_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_7127_)
);

FILL FILL_0__13484_ (
);

FILL FILL_0__13064_ (
);

FILL FILL380000x138320 (
);

FILL FILL282720x24700 (
);

FILL FILL257640x360620 (
);

OR2X2 _19419_ (
    .A(_8313_),
    .B(_8312_),
    .Y(_8314_)
);

FILL FILL_0__14689_ (
);

AND2X2 _14974_ (
    .A(_3995_),
    .B(_3994_),
    .Y(_3936_[29])
);

FILL FILL_0__14269_ (
);

AND2X2 _14554_ (
    .A(_3775_),
    .B(_3774_),
    .Y(_3738_[18])
);

OR2X2 _14134_ (
    .A(_3534_),
    .B(_3531_),
    .Y(\datapath_1.alu_1.ALUInB [30])
);

FILL FILL220400x103740 (
);

FILL FILL_0__15630_ (
);

FILL FILL_0__15210_ (
);

FILL FILL274360x276640 (
);

FILL FILL124640x34580 (
);

OR2X2 _15759_ (
    .A(_4708_),
    .B(_4707_),
    .Y(_4709_)
);

OR2X2 _15339_ (
    .A(_4294_),
    .B(_4295_),
    .Y(_4296_)
);

DFFSR _10894_ (
    .CLK(clk_bF$buf4),
    .D(_1191_[19]),
    .Q(\datapath_1.regfile_1.regOut[19] [19]),
    .R(rst_bF$buf20),
    .S(vdd)
);

OR2X2 _10474_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .B(_1058__bF$buf4),
    .Y(_1048_)
);

FILL FILL_1__17002_ (
);

OR2X2 _10054_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .B(_860__bF$buf4),
    .Y(_828_)
);

FILL FILL_0__16835_ (
);

AND2X2 _16700_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_5635_)
);

FILL FILL71440x4940 (
);

FILL FILL_0__11130_ (
);

OR2X2 _19172_ (
    .A(_8066_),
    .B(_8069_),
    .Y(_8070_)
);

FILL FILL490200x39520 (
);

OR2X2 _8622_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_93_)
);

FILL FILL_1__18627_ (
);

DFFSR _11679_ (
    .CLK(clk_bF$buf107),
    .D(_1587_[30]),
    .Q(\datapath_1.regfile_1.regOut[25] [30]),
    .R(rst_bF$buf56),
    .S(vdd)
);

OR2X2 _11259_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_1451_)
);

FILL FILL_1__13342_ (
);

AND2X2 _17905_ (
    .A(_6328__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_6823_)
);

AND2X2 _12620_ (
    .A(_2184_),
    .B(_2174_),
    .Y(_2185_)
);

AND2X2 _12200_ (
    .A(_1918_),
    .B(_1981_),
    .Y(_1917_[0])
);

AND2X2 _15092_ (
    .A(_4075_),
    .B(_4066_),
    .Y(_4076_)
);

FILL FILL128440x34580 (
);

FILL FILL171000x266760 (
);

AND2X2 _9827_ (
    .A(_716_),
    .B(_715_),
    .Y(_663_[26])
);

AND2X2 _9407_ (
    .A(_496_),
    .B(_495_),
    .Y(_465_[15])
);

FILL FILL249280x281580 (
);

FILL FILL255360x222300 (
);

FILL FILL_1__14547_ (
);

OR2X2 _13825_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [3]),
    .Y(_3283_)
);

FILL FILL437760x29640 (
);

AND2X2 _13405_ (
    .A(_2940_),
    .B(_2938_),
    .Y(_2941_)
);

AND2X2 _16297_ (
    .A(_4151__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_5239_)
);

FILL FILL310080x345800 (
);

FILL FILL_0__17373_ (
);

FILL FILL53200x187720 (
);

FILL FILL_1__10047_ (
);

OR2X2 _9580_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .B(_596__bF$buf3),
    .Y(_592_)
);

OR2X2 _9160_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .B(_398__bF$buf4),
    .Y(_372_)
);

FILL FILL67640x148200 (
);

FILL FILL_0__10821_ (
);

FILL FILL_0__10401_ (
);

FILL FILL266760x19760 (
);

FILL FILL_0__18578_ (
);

OR2X2 _18863_ (
    .A(_7765_),
    .B(_7764_),
    .Y(_7766_)
);

FILL FILL_0__18158_ (
);

FILL FILL_0_BUFX2_insert801 (
);

AND2X2 _18443_ (
    .A(_6206__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_7353_)
);

OR2X2 _18023_ (
    .A(_6931_),
    .B(_6938_),
    .Y(_6939_)
);

FILL FILL_0_BUFX2_insert803 (
);

FILL FILL_0__13293_ (
);

FILL FILL_0_BUFX2_insert805 (
);

FILL FILL_0_BUFX2_insert806 (
);

FILL FILL_0_BUFX2_insert807 (
);

FILL FILL_0_BUFX2_insert808 (
);

FILL FILL112480x103740 (
);

FILL FILL_0_BUFX2_insert809 (
);

FILL FILL_0__8679_ (
);

OR2X2 _19228_ (
    .A(_8093_),
    .B(_8125_),
    .Y(_8126_)
);

OR2X2 _14783_ (
    .A(vdd),
    .B(_2_[9]),
    .Y(_3888_)
);

FILL FILL_0__14498_ (
);

DFFSR _14363_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[27]),
    .Q(ALUOut[27]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL38760x232180 (
);

FILL FILL_1__13818_ (
);

FILL FILL38000x330980 (
);

FILL FILL370120x202540 (
);

FILL FILL314640x14820 (
);

AND2X2 _15988_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_4935_)
);

OR2X2 _15568_ (
    .A(_4517_),
    .B(_4520_),
    .Y(_4521_)
);

AND2X2 _15148_ (
    .A(_4114_),
    .B(_4016_),
    .Y(_4115_)
);

FILL FILL_1__17651_ (
);

FILL FILL_1__17231_ (
);

AND2X2 _10283_ (
    .A(_940_),
    .B(_939_),
    .Y(_927_[6])
);

FILL FILL107160x14820 (
);

FILL FILL501600x79040 (
);

FILL FILL_0__16224_ (
);

FILL FILL177840x108680 (
);

FILL FILL81320x281580 (
);

OR2X2 _8851_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .B(_266__bF$buf0),
    .Y(_206_)
);

BUFX2 _8431_ (
    .A(_2_[7]),
    .Y(memoryWriteData[7])
);

OR2X2 _11488_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .B(_1586__bF$buf0),
    .Y(_1564_)
);

OR2X2 _11068_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .B(_1388__bF$buf1),
    .Y(_1344_)
);

FILL FILL_1__13991_ (
);

FILL FILL_0__17849_ (
);

FILL FILL_0__17429_ (
);

OR2X2 _17714_ (
    .A(_6634_),
    .B(_6633_),
    .Y(_6635_)
);

FILL FILL_0__12564_ (
);

FILL FILL_0__12144_ (
);

OR2X2 _9636_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_609_)
);

DFFSR _9216_ (
    .CLK(clk_bF$buf106),
    .D(_333_[18]),
    .Q(\datapath_1.regfile_1.regOut[6] [18]),
    .R(rst_bF$buf96),
    .S(vdd)
);

FILL FILL299440x247000 (
);

FILL FILL59280x256880 (
);

OR2X2 _18919_ (
    .A(_7820_),
    .B(_7817_),
    .Y(_7821_)
);

FILL FILL228760x49400 (
);

FILL FILL_0__13769_ (
);

FILL FILL_0__13349_ (
);

AND2X2 _13634_ (
    .A(_3084__bF$buf3),
    .B(\aluControl_1.inst [4]),
    .Y(_3123_)
);

NOR3X1 _13214_ (
    .A(_2761_),
    .B(_2757_),
    .C(_2759_),
    .Y(_2762_)
);

FILL FILL285760x271700 (
);

FILL FILL_0__14710_ (
);

FILL FILL448400x232180 (
);

FILL FILL_1__9798_ (
);

FILL FILL311600x266760 (
);

FILL FILL_0__17182_ (
);

FILL FILL308560x217360 (
);

AND2X2 _14839_ (
    .A(_3925_),
    .B(_3924_),
    .Y(_3870_[27])
);

AND2X2 _14419_ (
    .A(_3705_),
    .B(_3704_),
    .Y(_3672_[16])
);

FILL FILL_0__15915_ (
);

FILL FILL167200x19760 (
);

FILL FILL_0__10210_ (
);

OR2X2 _18672_ (
    .A(_7577_),
    .B(_7576_),
    .Y(_7578_)
);

OR2X2 _18252_ (
    .A(_7148_),
    .B(_7164_),
    .Y(_7165_)
);

FILL FILL_0__8488_ (
);

DFFSR _10759_ (
    .CLK(clk_bF$buf47),
    .D(_1125_[13]),
    .Q(\datapath_1.regfile_1.regOut[18] [13]),
    .R(rst_bF$buf51),
    .S(vdd)
);

OR2X2 _10339_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .B(_992__bF$buf2),
    .Y(_978_)
);

FILL FILL_1__12842_ (
);

FILL FILL_1__12422_ (
);

FILL FILL_0__11835_ (
);

OR2X2 _11700_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_1665_)
);

OR2X2 _19457_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_8340_)
);

AND2X2 _19037_ (
    .A(_6302__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_7937_)
);

OR2X2 _14592_ (
    .A(memoryOutData[31]),
    .B(_3803__bF$buf1),
    .Y(_3801_)
);

AND2X2 _14172_ (
    .A(_3559_),
    .B(_3558_),
    .Y(\datapath_1.mux_wd3.dout [9])
);

OR2X2 _8907_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_243_)
);

FILL FILL70680x207480 (
);

FILL FILL364800x172900 (
);

FILL FILL_1__13207_ (
);

FILL FILL374680x118560 (
);

OR2X2 _12905_ (
    .A(_2469_),
    .B(_2450_),
    .Y(_2470_)
);

FILL FILL_1_BUFX2_insert358 (
);

OR2X2 _15797_ (
    .A(_4745_),
    .B(_4746_),
    .Y(_4747_)
);

AND2X2 _15377_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_4333_)
);

FILL FILL_1__17880_ (
);

OR2X2 _10092_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_853_)
);

FILL FILL148200x158080 (
);

FILL FILL125400x49400 (
);

FILL FILL_0__16873_ (
);

FILL FILL_0__16453_ (
);

FILL FILL_0__16033_ (
);

FILL FILL55480x286520 (
);

AND2X2 _8660_ (
    .A(_118_),
    .B(_117_),
    .Y(_69_[24])
);

AND2X2 _11297_ (
    .A(_1456_),
    .B(_1519_),
    .Y(_1455_[0])
);

OR2X2 _17943_ (
    .A(_6858_),
    .B(_6859_),
    .Y(_6860_)
);

FILL FILL_0__17658_ (
);

FILL FILL_0__17238_ (
);

AND2X2 _17523_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_6447_)
);

OR2X2 _17103_ (
    .A(_6030_),
    .B(_6031_),
    .Y(_6032_)
);

FILL FILL_0__12793_ (
);

FILL FILL_0__12373_ (
);

FILL FILL313120x370500 (
);

FILL FILL427120x118560 (
);

DFFSR _9865_ (
    .CLK(clk_bF$buf74),
    .D(_663_[22]),
    .Q(\datapath_1.regfile_1.regOut[11] [22]),
    .R(rst_bF$buf47),
    .S(vdd)
);

OR2X2 _9445_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .B(_530__bF$buf0),
    .Y(_522_)
);

OR2X2 _9025_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .B(_332__bF$buf0),
    .Y(_302_)
);

FILL FILL203680x266760 (
);

FILL FILL_1__14165_ (
);

FILL FILL129200x49400 (
);

AND2X2 _18728_ (
    .A(_6211__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_7633_)
);

OR2X2 _18308_ (
    .A(_7219_),
    .B(_7216_),
    .Y(_7220_)
);

FILL FILL_0__13998_ (
);

AND2X2 _13863_ (
    .A(_3308_),
    .B(_3307_),
    .Y(\datapath_1.alu_1.ALUInA [15])
);

FILL FILL_0__13158_ (
);

AND2X2 _13443_ (
    .A(_2634_),
    .B(_2752_),
    .Y(_2976_)
);

OAI21X1 _13023_ (
    .A(_2332_),
    .B(\datapath_1.alu_1.ALUInB [24]),
    .C(_2476_),
    .Y(_2582_)
);

FILL FILL52440x182780 (
);

FILL FILL80560x54340 (
);

FILL FILL_0__9905_ (
);

FILL FILL34960x355680 (
);

FILL FILL256120x187720 (
);

OR2X2 _14648_ (
    .A(vdd),
    .B(\datapath_1.a [7]),
    .Y(_3818_)
);

OR2X2 _14228_ (
    .A(\datapath_1.Data [28]),
    .B(_3605__bF$buf3),
    .Y(_3597_)
);

FILL FILL_1__16731_ (
);

FILL FILL_0__15724_ (
);

FILL FILL_0__15304_ (
);

FILL FILL273600x197600 (
);

FILL FILL_0__18196_ (
);

AND2X2 _18481_ (
    .A(_6282__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_7390_)
);

AND2X2 _18061_ (
    .A(_6244__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_6976_)
);

FILL FILL100320x256880 (
);

AND2X2 _10988_ (
    .A(_1310_),
    .B(_1309_),
    .Y(_1257_[26])
);

AND2X2 _10568_ (
    .A(_1090_),
    .B(_1089_),
    .Y(_1059_[15])
);

AND2X2 _10148_ (
    .A(_870_),
    .B(_869_),
    .Y(_861_[4])
);

FILL FILL_1__12231_ (
);

FILL FILL_0__16929_ (
);

FILL FILL_0__11644_ (
);

FILL FILL_0__11224_ (
);

AND2X2 _19266_ (
    .A(_6317__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_8163_)
);

FILL FILL127680x163020 (
);

OR2X2 _8716_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_200__bF$buf0),
    .Y(_136_)
);

FILL FILL161880x4940 (
);

FILL FILL371640x49400 (
);

FILL FILL488680x138320 (
);

FILL FILL9880x261820 (
);

FILL FILL_1__13856_ (
);

OR2X2 _12714_ (
    .A(\datapath_1.alu_1.ALUInA [19]),
    .B(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2279_)
);

FILL FILL85880x0 (
);

FILL FILL442320x311220 (
);

INVX1 _15186_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .Y(_4144_)
);

FILL FILL319960x212420 (
);

FILL FILL_1_BUFX2_insert27 (
);

FILL FILL_1_BUFX2_insert29 (
);

FILL FILL291840x64220 (
);

FILL FILL_0__16682_ (
);

FILL FILL22800x271700 (
);

FILL FILL429400x98800 (
);

NOR2X1 _13919_ (
    .A(ALUSrcB[0]),
    .B(ALUSrcB[1]),
    .Y(_3350_)
);

FILL FILL466640x74100 (
);

FILL FILL_1__18054_ (
);

FILL FILL_0__17887_ (
);

AND2X2 _17752_ (
    .A(_6262__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_6672_)
);

FILL FILL_0__17047_ (
);

NOR2X1 _17332_ (
    .A(_6257_),
    .B(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_6258_)
);

AND2X2 _9674_ (
    .A(_634_),
    .B(_633_),
    .Y(_597_[18])
);

AND2X2 _9254_ (
    .A(_414_),
    .B(_413_),
    .Y(_399_[7])
);

FILL FILL_1__11502_ (
);

FILL FILL_0__10915_ (
);

OR2X2 _18957_ (
    .A(_7858_),
    .B(_7856_),
    .Y(_7859_)
);

AND2X2 _18537_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_7445_)
);

AND2X2 _18117_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_7032_)
);

FILL FILL_0__13387_ (
);

AND2X2 _13672_ (
    .A(_3089__bF$buf1),
    .B(gnd),
    .Y(_3156_)
);

NOR2X1 _13252_ (
    .A(_2435_),
    .B(_2498_),
    .Y(_2797_)
);

FILL FILL_1_BUFX2_insert1117 (
);

FILL FILL_1_BUFX2_insert1119 (
);

FILL FILL_1__12707_ (
);

FILL FILL303240x113620 (
);

FILL FILL328320x158080 (
);

FILL FILL415720x163020 (
);

FILL FILL85880x123500 (
);

DFFSR _14877_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[25]),
    .Q(_2_[25]),
    .R(rst_bF$buf61),
    .S(vdd)
);

OR2X2 _14457_ (
    .A(memoryOutData[29]),
    .B(_3737__bF$buf0),
    .Y(_3731_)
);

AND2X2 _14037_ (
    .A(_3344__bF$buf2),
    .B(gnd),
    .Y(_3451_)
);

FILL FILL480320x345800 (
);

FILL FILL_1__16120_ (
);

FILL FILL_0__15953_ (
);

AND2X2 _18290_ (
    .A(_6255__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_7202_)
);

FILL FILL44840x19760 (
);

FILL FILL329080x34580 (
);

FILL FILL142880x222300 (
);

FILL FILL_1__17745_ (
);

OR2X2 _10797_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_1203_)
);

DFFSR _10377_ (
    .CLK(clk_bF$buf61),
    .D(_927_[18]),
    .Q(\datapath_1.regfile_1.regOut[15] [18]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL250040x355680 (
);

FILL FILL_0__16738_ (
);

FILL FILL438520x113620 (
);

AND2X2 _16603_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_5540_)
);

FILL FILL_0__16318_ (
);

FILL FILL_0__11873_ (
);

FILL FILL_0__11453_ (
);

AND2X2 _19495_ (
    .A(_8365_),
    .B(_8364_),
    .Y(_8320_[22])
);

AND2X2 _19075_ (
    .A(_6315__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_7975_)
);

DFFSR _8945_ (
    .CLK(clk_bF$buf59),
    .D(_201_[5]),
    .Q(\datapath_1.regfile_1.regOut[4] [5]),
    .R(rst_bF$buf106),
    .S(vdd)
);

AND2X2 _8525_ (
    .A(_48_),
    .B(_47_),
    .Y(_3_[22])
);

FILL FILL45600x365560 (
);

OR2X2 _17808_ (
    .A(_6722_),
    .B(_6726_),
    .Y(_6727_)
);

FILL FILL_0__12658_ (
);

NOR3X1 _12943_ (
    .A(_2506_),
    .B(_2499_),
    .C(_2502_),
    .Y(_2507_)
);

FILL FILL301720x44460 (
);

FILL FILL_0__12238_ (
);

INVX1 _12523_ (
    .A(\control_1.op [0]),
    .Y(_2113_)
);

OR2X2 _12103_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .B(_1916__bF$buf0),
    .Y(_1874_)
);

FILL FILL_1_BUFX2_insert737 (
);

FILL FILL350360x172900 (
);

FILL FILL_1_BUFX2_insert739 (
);

FILL FILL436240x187720 (
);

FILL FILL_0__16491_ (
);

FILL FILL_0__16071_ (
);

AND2X2 _13728_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3204_)
);

FILL FILL206720x291460 (
);

FILL FILL162640x9880 (
);

OAI21X1 _13308_ (
    .A(_2172_),
    .B(_2171_),
    .C(_2169_),
    .Y(_2849_)
);

BUFX2 BUFX2_insert400 (
    .A(_6297_),
    .Y(_6297__bF$buf0)
);

BUFX2 BUFX2_insert401 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf4 )
);

BUFX2 BUFX2_insert402 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf3 )
);

BUFX2 BUFX2_insert403 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf2 )
);

BUFX2 BUFX2_insert404 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf1 )
);

AND2X2 _17981_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_6898_)
);

FILL FILL_0__17696_ (
);

AND2X2 _17561_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_6484_)
);

BUFX2 BUFX2_insert405 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf0 )
);

FILL FILL_0__17276_ (
);

BUFX2 BUFX2_insert406 (
    .A(_4172_),
    .Y(_4172__bF$buf4)
);

OR2X2 _17141_ (
    .A(_6069_),
    .B(_6068_),
    .Y(_6070_)
);

BUFX2 BUFX2_insert407 (
    .A(_4172_),
    .Y(_4172__bF$buf3)
);

BUFX2 BUFX2_insert408 (
    .A(_4172_),
    .Y(_4172__bF$buf2)
);

BUFX2 BUFX2_insert409 (
    .A(_4172_),
    .Y(_4172__bF$buf1)
);

DFFSR _9483_ (
    .CLK(clk_bF$buf66),
    .D(_465_[27]),
    .Q(\datapath_1.regfile_1.regOut[8] [27]),
    .R(rst_bF$buf80),
    .S(vdd)
);

OR2X2 _9063_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_327_)
);

FILL FILL279680x59280 (
);

FILL FILL_1__11311_ (
);

FILL FILL_1__19068_ (
);

FILL FILL_0__10724_ (
);

OR2X2 _18766_ (
    .A(_7669_),
    .B(_7670_),
    .Y(_7671_)
);

FILL FILL500080x123500 (
);

AND2X2 _18346_ (
    .A(_6236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_7257_)
);

FILL FILL232560x29640 (
);

AND2X2 _13481_ (
    .A(_3010_),
    .B(_3009_),
    .Y(\datapath_1.a3 [2])
);

OR2X2 _13061_ (
    .A(_2613_),
    .B(_2617_),
    .Y(_2618_)
);

FILL FILL_0__19002_ (
);

FILL FILL164920x4940 (
);

FILL FILL_1__12936_ (
);

FILL FILL261440x123500 (
);

FILL FILL407360x39520 (
);

FILL FILL_0__9943_ (
);

FILL FILL_0__9523_ (
);

FILL FILL_0__11509_ (
);

FILL FILL_0__9103_ (
);

FILL FILL60800x237120 (
);

AND2X2 _14686_ (
    .A(_3843_),
    .B(_3842_),
    .Y(_3804_[19])
);

AND2X2 _14266_ (
    .A(_3623_),
    .B(_3622_),
    .Y(_3606_[8])
);

FILL FILL117800x242060 (
);

FILL FILL_0__15342_ (
);

FILL FILL32680x0 (
);

OR2X2 _10186_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_926__bF$buf0),
    .Y(_896_)
);

FILL FILL_0__16967_ (
);

FILL FILL_0__16547_ (
);

OR2X2 _16832_ (
    .A(_5763_),
    .B(_5764_),
    .Y(_5765_)
);

OR2X2 _16412_ (
    .A(_5351_),
    .B(_5350_),
    .Y(_5352_)
);

FILL FILL_0__16127_ (
);

FILL FILL117800x108680 (
);

FILL FILL104120x247000 (
);

FILL FILL47120x335920 (
);

FILL FILL_0__11682_ (
);

FILL FILL18240x232180 (
);

OR2X2 _8754_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_161_)
);

FILL FILL383800x59280 (
);

FILL FILL235600x326040 (
);

NOR2X1 _17617_ (
    .A(_6310__bF$buf1),
    .B(_6538_),
    .Y(_6539_)
);

FILL FILL422560x143260 (
);

FILL FILL_0__12887_ (
);

FILL FILL166440x133380 (
);

AND2X2 _12752_ (
    .A(_2287_),
    .B(_2316_),
    .Y(_2317_)
);

AND2X2 _12332_ (
    .A(_1986_),
    .B(_1985_),
    .Y(_1983_[1])
);

FILL FILL394440x197600 (
);

AND2X2 _9959_ (
    .A(_784_),
    .B(_783_),
    .Y(_729_[27])
);

FILL FILL322240x237120 (
);

AND2X2 _9539_ (
    .A(_564_),
    .B(_563_),
    .Y(_531_[16])
);

AND2X2 _9119_ (
    .A(_344_),
    .B(_343_),
    .Y(_333_[5])
);

FILL FILL_1__8496_ (
);

FILL FILL202920x187720 (
);

FILL FILL183920x143260 (
);

FILL FILL221160x256880 (
);

FILL FILL239400x247000 (
);

FILL FILL_1__14259_ (
);

FILL FILL_0_BUFX2_insert390 (
);

FILL FILL_0_BUFX2_insert391 (
);

FILL FILL_0_BUFX2_insert392 (
);

FILL FILL35720x108680 (
);

AND2X2 _13957_ (
    .A(_3352__bF$buf1),
    .B(\aluControl_1.inst [3]),
    .Y(_3383_)
);

FILL FILL_0_BUFX2_insert394 (
);

OR2X2 _13537_ (
    .A(IorD_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [16]),
    .Y(_3046_)
);

XOR2X1 _13117_ (
    .A(_2281_),
    .B(_2669_),
    .Y(_2670_)
);

FILL FILL_0_BUFX2_insert396 (
);

FILL FILL_0_BUFX2_insert398 (
);

FILL FILL_1__15200_ (
);

FILL FILL_1__18092_ (
);

AND2X2 _17790_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_6710_)
);

AND2X2 _17370_ (
    .A(_6295_),
    .B(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_6296_)
);

FILL FILL_1__10179_ (
);

FILL FILL426360x251940 (
);

OR2X2 _9292_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .B(_464__bF$buf3),
    .Y(_440_)
);

FILL FILL_0__15818_ (
);

FILL FILL_0__10953_ (
);

FILL FILL_0__10533_ (
);

FILL FILL443840x261820 (
);

AND2X2 _18995_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_7896_)
);

OR2X2 _18575_ (
    .A(_7479_),
    .B(_7482_),
    .Y(_7483_)
);

AND2X2 _18155_ (
    .A(_6282__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_7069_)
);

OAI21X1 _13290_ (
    .A(_2830_),
    .B(_2829_),
    .C(_2832_),
    .Y(_2833_)
);

FILL FILL148200x0 (
);

FILL FILL493240x316160 (
);

FILL FILL_0__19231_ (
);

FILL FILL_0__9752_ (
);

FILL FILL_0__11318_ (
);

AND2X2 _11603_ (
    .A(_1620_),
    .B(_1619_),
    .Y(_1587_[16])
);

FILL FILL73720x276640 (
);

DFFSR _14495_ (
    .CLK(clk_bF$buf20),
    .D(_3672_[30]),
    .Q(\datapath_1.Data [30]),
    .R(rst_bF$buf22),
    .S(vdd)
);

AND2X2 _14075_ (
    .A(_3350__bF$buf4),
    .B(_2_[22]),
    .Y(_3484_)
);

FILL FILL228000x54340 (
);

FILL FILL_0__15991_ (
);

FILL FILL145160x153140 (
);

FILL FILL_0__15571_ (
);

FILL FILL_0__15151_ (
);

FILL FILL200640x370500 (
);

OR2X2 _12808_ (
    .A(_2157__bF$buf0),
    .B(_2372_),
    .Y(_2373_)
);

FILL FILL_0__16776_ (
);

OR2X2 _16641_ (
    .A(_5573_),
    .B(_5576_),
    .Y(_5577_)
);

FILL FILL_0__16356_ (
);

AND2X2 _16221_ (
    .A(_4230__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_5164_)
);

FILL FILL_0__11071_ (
);

FILL FILL_1__9913_ (
);

OR2X2 _8983_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .B(_332__bF$buf4),
    .Y(_274_)
);

DFFSR _8563_ (
    .CLK(clk_bF$buf0),
    .D(_3_[10]),
    .Q(\datapath_1.regfile_1.regOut[1] [10]),
    .R(rst_bF$buf64),
    .S(vdd)
);

FILL FILL112480x98800 (
);

FILL FILL368600x0 (
);

FILL FILL346560x24700 (
);

FILL FILL_1__18568_ (
);

FILL FILL504640x375440 (
);

FILL FILL_1__13283_ (
);

FILL FILL435480x182780 (
);

FILL FILL380760x153140 (
);

OR2X2 _17846_ (
    .A(_6757_),
    .B(_6764_),
    .Y(_6765_)
);

AND2X2 _17426_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_6351_)
);

OR2X2 _17006_ (
    .A(_5935_),
    .B(_5936_),
    .Y(_5937_)
);

AND2X2 _12981_ (
    .A(_2541_),
    .B(_2342_),
    .Y(_2542_)
);

FILL FILL_0__12276_ (
);

AND2X2 _12561_ (
    .A(_2132_),
    .B(\control_1.op [2]),
    .Y(_2082_)
);

OR2X2 _12141_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_1899_)
);

FILL FILL_0__18502_ (
);

OR2X2 _9768_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_677_)
);

DFFSR _9348_ (
    .CLK(clk_bF$buf93),
    .D(_399_[21]),
    .Q(\datapath_1.regfile_1.regOut[7] [21]),
    .R(rst_bF$buf41),
    .S(vdd)
);

FILL FILL_0__8603_ (
);

AND2X2 _13766_ (
    .A(_3081__bF$buf2),
    .B(ALUOut[25]),
    .Y(_3236_)
);

NAND2X1 _13346_ (
    .A(_2187_),
    .B(_2873_),
    .Y(_2886_)
);

FILL FILL269800x296400 (
);

FILL FILL_0__14842_ (
);

FILL FILL_0__14422_ (
);

FILL FILL183160x187720 (
);

FILL FILL_0__9808_ (
);

FILL FILL37240x74100 (
);

FILL FILL_1__16214_ (
);

OR2X2 _15912_ (
    .A(_4852_),
    .B(_4859_),
    .Y(_4860_)
);

FILL FILL_0__15207_ (
);

FILL FILL_0__10342_ (
);

FILL FILL12160x311220 (
);

FILL FILL_0__18099_ (
);

OR2X2 _18384_ (
    .A(_7261_),
    .B(_7294_),
    .Y(_7295_)
);

FILL FILL159600x316160 (
);

FILL FILL_0__19460_ (
);

FILL FILL_0__19040_ (
);

FILL FILL474240x54340 (
);

FILL FILL_1__17419_ (
);

FILL FILL_1__12974_ (
);

FILL FILL_1__12554_ (
);

FILL FILL182400x83980 (
);

FILL FILL_0__11967_ (
);

FILL FILL_0__9141_ (
);

OR2X2 _11832_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_1733_)
);

DFFSR _11412_ (
    .CLK(clk_bF$buf21),
    .D(_1455_[21]),
    .Q(\datapath_1.regfile_1.regOut[23] [21]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL456000x103740 (
);

AND2X2 _19169_ (
    .A(_6271__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_8067_)
);

FILL FILL171760x281580 (
);

OR2X2 _8619_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_91_)
);

FILL FILL357200x93860 (
);

XOR2X1 _12617_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2182_)
);

AND2X2 _15089_ (
    .A(_4029_),
    .B(_4041_),
    .Y(_4074_)
);

FILL FILL_1__17172_ (
);

OR2X2 _16870_ (
    .A(_5802_),
    .B(_5801_),
    .Y(_5803_)
);

FILL FILL_0__16165_ (
);

AND2X2 _16450_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_5389_)
);

AND2X2 _16030_ (
    .A(_4167__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_4976_)
);

FILL FILL_1__9302_ (
);

AND2X2 _8792_ (
    .A(_186_),
    .B(_185_),
    .Y(_135_[25])
);

FILL FILL224200x281580 (
);

FILL FILL_1__10200_ (
);

FILL FILL267520x345800 (
);

AND2X2 _17655_ (
    .A(_6289__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_6577_)
);

OR2X2 _17235_ (
    .A(_6160_),
    .B(_6161_),
    .Y(_6162_)
);

INVX1 _12790_ (
    .A(_2354_),
    .Y(_2355_)
);

OR2X2 _12370_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .B(_2048__bF$buf3),
    .Y(_2012_)
);

FILL FILL_0__12085_ (
);

FILL FILL238640x242060 (
);

FILL FILL_0__18731_ (
);

FILL FILL_0__18311_ (
);

DFFSR _9997_ (
    .CLK(clk_bF$buf93),
    .D(_729_[25]),
    .Q(\datapath_1.regfile_1.regOut[12] [25]),
    .R(rst_bF$buf41),
    .S(vdd)
);

OR2X2 _9577_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .B(_596__bF$buf4),
    .Y(_590_)
);

OR2X2 _9157_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .B(_398__bF$buf2),
    .Y(_370_)
);

FILL FILL107160x350740 (
);

FILL FILL_0__8412_ (
);

FILL FILL_1__14297_ (
);

FILL FILL_0_BUFX2_insert770 (
);

FILL FILL_0_BUFX2_insert771 (
);

FILL FILL_0_BUFX2_insert772 (
);

FILL FILL_0_BUFX2_insert774 (
);

AND2X2 _13995_ (
    .A(_3344__bF$buf3),
    .B(gnd),
    .Y(_3415_)
);

AND2X2 _13575_ (
    .A(_3071_),
    .B(_3070_),
    .Y(_1_[28])
);

NOR3X1 _13155_ (
    .A(_2702_),
    .B(_2703_),
    .C(_2705_),
    .Y(_2706_)
);

FILL FILL_0_BUFX2_insert776 (
);

FILL FILL_0_BUFX2_insert778 (
);

FILL FILL_0__19516_ (
);

FILL FILL_0__14231_ (
);

FILL FILL_0__9617_ (
);

FILL FILL_1__16863_ (
);

FILL FILL_0__15856_ (
);

FILL FILL_0__15436_ (
);

AND2X2 _15721_ (
    .A(_4135__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_4672_)
);

FILL FILL_0__15016_ (
);

AND2X2 _15301_ (
    .A(_4214__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_4258_)
);

FILL FILL_0__10571_ (
);

FILL FILL_0__10151_ (
);

OR2X2 _18193_ (
    .A(_7105_),
    .B(_7104_),
    .Y(_7106_)
);

FILL FILL_1__12363_ (
);

AND2X2 _16926_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_5858_)
);

AND2X2 _16506_ (
    .A(_5444_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd2 [19])
);

FILL FILL_0__9790_ (
);

FILL FILL_0__11776_ (
);

FILL FILL_0__11356_ (
);

OR2X2 _11641_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .B(_1652__bF$buf4),
    .Y(_1646_)
);

OR2X2 _11221_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_1454__bF$buf0),
    .Y(_1426_)
);

OR2X2 _19398_ (
    .A(_8292_),
    .B(_8289_),
    .Y(_8293_)
);

OR2X2 _8848_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_266__bF$buf2),
    .Y(_204_)
);

BUFX2 _8428_ (
    .A(_2_[4]),
    .Y(memoryWriteData[4])
);

FILL FILL276640x276640 (
);

FILL FILL147440x34580 (
);

FILL FILL_1__13148_ (
);

OR2X2 _12846_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2411_)
);

DFFSR _12426_ (
    .CLK(clk_bF$buf44),
    .D(_1983_[3]),
    .Q(\datapath_1.regfile_1.regOut[31] [3]),
    .R(rst_bF$buf16),
    .S(vdd)
);

OR2X2 _12006_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_1829_)
);

FILL FILL53200x232180 (
);

FILL FILL_0__13922_ (
);

FILL FILL_0__16394_ (
);

FILL FILL_1__9111_ (
);

FILL FILL422560x306280 (
);

FILL FILL_1__15714_ (
);

FILL FILL339720x316160 (
);

FILL FILL_0__14707_ (
);

FILL FILL_1__18186_ (
);

AND2X2 _17884_ (
    .A(_6312__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_6802_)
);

AND2X2 _17464_ (
    .A(_6302__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_6389_)
);

FILL FILL_0__17179_ (
);

AND2X2 _17044_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_5974_)
);

FILL FILL_0__18960_ (
);

FILL FILL_0__18540_ (
);

FILL FILL_0__18120_ (
);

FILL FILL257640x222300 (
);

AND2X2 _9386_ (
    .A(_482_),
    .B(_481_),
    .Y(_465_[8])
);

FILL FILL_1__11634_ (
);

OR2X2 _10912_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_1322__bF$buf0),
    .Y(_1260_)
);

FILL FILL_0__10207_ (
);

OR2X2 _18669_ (
    .A(_7574_),
    .B(_7573_),
    .Y(_7575_)
);

OR2X2 _18249_ (
    .A(_7160_),
    .B(_7161_),
    .Y(_7162_)
);

XOR2X1 _13384_ (
    .A(_2393_),
    .B(_2920_),
    .Y(_2921_)
);

FILL FILL_0__13099_ (
);

FILL FILL_0__19325_ (
);

FILL FILL_0__14460_ (
);

FILL FILL_0__14040_ (
);

FILL FILL391400x256880 (
);

FILL FILL_0__9426_ (
);

FILL FILL465120x172900 (
);

FILL FILL212800x192660 (
);

OR2X2 _14589_ (
    .A(memoryOutData[30]),
    .B(_3803__bF$buf1),
    .Y(_3799_)
);

AND2X2 _14169_ (
    .A(_3557_),
    .B(_3556_),
    .Y(\datapath_1.mux_wd3.dout [8])
);

FILL FILL459040x9880 (
);

FILL FILL_1__16672_ (
);

AND2X2 _15950_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_4897_)
);

FILL FILL_0__15665_ (
);

AND2X2 _15530_ (
    .A(_4183__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_4484_)
);

FILL FILL_0__15245_ (
);

NAND3X1 _15110_ (
    .A(_4013_),
    .B(_4054_),
    .C(_4017_),
    .Y(_4090_)
);

FILL FILL23560x93860 (
);

FILL FILL424080x83980 (
);

FILL FILL_1__17037_ (
);

OR2X2 _10089_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_851_)
);

FILL FILL262960x9880 (
);

OR2X2 _16735_ (
    .A(_5668_),
    .B(_5669_),
    .Y(_5670_)
);

AND2X2 _16315_ (
    .A(_4187__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_5256_)
);

AND2X2 _11870_ (
    .A(_1758_),
    .B(_1757_),
    .Y(_1719_[19])
);

FILL FILL_0__11585_ (
);

AND2X2 _11450_ (
    .A(_1538_),
    .B(_1537_),
    .Y(_1521_[8])
);

DFFSR _11030_ (
    .CLK(clk_bF$buf55),
    .D(_1257_[26]),
    .Q(\datapath_1.regfile_1.regOut[20] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

FILL FILL427880x133380 (
);

FILL FILL_0__17811_ (
);

FILL FILL262960x0 (
);

AND2X2 _8657_ (
    .A(_116_),
    .B(_115_),
    .Y(_69_[23])
);

FILL FILL112480x177840 (
);

FILL FILL372400x202540 (
);

FILL FILL_1__13797_ (
);

FILL FILL_1__13377_ (
);

NAND2X1 _12655_ (
    .A(_2218_),
    .B(_2219_),
    .Y(_2220_)
);

OR2X2 _12235_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .B(_1982__bF$buf0),
    .Y(_1942_)
);

FILL FILL_0__13311_ (
);

FILL FILL376200x123500 (
);

FILL FILL_0_BUFX2_insert1121 (
);

FILL FILL_0_BUFX2_insert1123 (
);

FILL FILL_0_BUFX2_insert1124 (
);

FILL FILL_0_BUFX2_insert1125 (
);

FILL FILL_0_BUFX2_insert1126 (
);

FILL FILL_0_BUFX2_insert1127 (
);

FILL FILL_0_BUFX2_insert1129 (
);

FILL FILL297920x326040 (
);

OR2X2 _14801_ (
    .A(vdd),
    .B(_2_[15]),
    .Y(_3900_)
);

FILL FILL_0__14516_ (
);

AND2X2 _17693_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_6614_)
);

OR2X2 _17273_ (
    .A(_6199_),
    .B(_6168_),
    .Y(_6200_)
);

FILL FILL201400x350740 (
);

OR2X2 _9195_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_395_)
);

FILL FILL_1__11443_ (
);

FILL FILL_0__10856_ (
);

AND2X2 _10721_ (
    .A(_1172_),
    .B(_1171_),
    .Y(_1125_[23])
);

FILL FILL_0__10016_ (
);

AND2X2 _10301_ (
    .A(_952_),
    .B(_951_),
    .Y(_927_[12])
);

AND2X2 _18898_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_7801_)
);

OR2X2 _18478_ (
    .A(_7383_),
    .B(_7386_),
    .Y(_7387_)
);

OR2X2 _18058_ (
    .A(_6941_),
    .B(_6973_),
    .Y(_6974_)
);

NAND2X1 _13193_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2742_)
);

FILL FILL224960x202540 (
);

FILL FILL64600x54340 (
);

FILL FILL_0__9655_ (
);

FILL FILL_0__9235_ (
);

DFFSR _11926_ (
    .CLK(clk_bF$buf69),
    .D(_1719_[19]),
    .Q(\datapath_1.regfile_1.regOut[27] [19]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL505400x355680 (
);

OR2X2 _11506_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_1586__bF$buf1),
    .Y(_1576_)
);

FILL FILL345040x281580 (
);

FILL FILL85880x93860 (
);

FILL FILL351120x222300 (
);

FILL FILL381520x133380 (
);

AND2X2 _14398_ (
    .A(_3691_),
    .B(_3690_),
    .Y(_3672_[9])
);

FILL FILL437000x237120 (
);

FILL FILL_0__15894_ (
);

FILL FILL241680x118560 (
);

FILL FILL_0__15474_ (
);

FILL FILL281200x227240 (
);

FILL FILL_1__8611_ (
);

FILL FILL139840x286520 (
);

FILL FILL_1__17686_ (
);

FILL FILL158080x355680 (
);

OR2X2 _16964_ (
    .A(_5893_),
    .B(_5894_),
    .Y(_5895_)
);

OR2X2 _16544_ (
    .A(_5478_),
    .B(_5481_),
    .Y(_5482_)
);

FILL FILL_0__16259_ (
);

AND2X2 _16124_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_5068_)
);

FILL FILL81320x330980 (
);

FILL FILL_0__17620_ (
);

FILL FILL_0__17200_ (
);

FILL FILL72960x207480 (
);

OR2X2 _8886_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_229_)
);

OR2X2 _8466_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_9_)
);

FILL FILL89680x93860 (
);

FILL FILL376960x118560 (
);

OR2X2 _17749_ (
    .A(_6667_),
    .B(_6668_),
    .Y(_6669_)
);

AND2X2 _17329_ (
    .A(_6254_),
    .B(_6201_),
    .Y(_6255_)
);

FILL FILL_0__12599_ (
);

AND2X2 _12884_ (
    .A(_2430_),
    .B(_2448_),
    .Y(_2449_)
);

NOR2X1 _12464_ (
    .A(_2057_),
    .B(_2052_),
    .Y(ALUControl[0])
);

DFFSR _12044_ (
    .CLK(clk_bF$buf67),
    .D(_1785_[8]),
    .Q(\datapath_1.regfile_1.regOut[28] [8]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL_0__18825_ (
);

FILL FILL_0__18405_ (
);

FILL FILL_0__13960_ (
);

FILL FILL_0__13540_ (
);

FILL FILL311600x128440 (
);

FILL FILL_0__8926_ (
);

FILL FILL_0__8506_ (
);

FILL FILL_1_BUFX2_insert1080 (
);

FILL FILL_1_BUFX2_insert1082 (
);

FILL FILL_1_BUFX2_insert1084 (
);

AND2X2 _13669_ (
    .A(_3084__bF$buf3),
    .B(\datapath_1.PCJump [11]),
    .Y(_3153_)
);

XOR2X1 _13249_ (
    .A(_2235_),
    .B(_2793_),
    .Y(_2794_)
);

FILL FILL_1__15332_ (
);

DFFSR _14610_ (
    .CLK(clk_bF$buf31),
    .D(_3738_[16]),
    .Q(\datapath_1.PCJump [18]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _17082_ (
    .A(_6011_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [28])
);

FILL FILL_1__16537_ (
);

FILL FILL_1__11252_ (
);

OR2X2 _15815_ (
    .A(_4763_),
    .B(_4762_),
    .Y(_4764_)
);

OR2X2 _10950_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_1285_)
);

FILL FILL_0__10665_ (
);

OR2X2 _10530_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_1065_)
);

FILL FILL54720x182780 (
);

DFFSR _10110_ (
    .CLK(clk_bF$buf75),
    .D(_795_[9]),
    .Q(\datapath_1.regfile_1.regOut[13] [9]),
    .R(rst_bF$buf24),
    .S(vdd)
);

AND2X2 _18287_ (
    .A(_6259__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_7199_)
);

FILL FILL478040x143260 (
);

FILL FILL383040x103740 (
);

FILL FILL258400x187720 (
);

FILL FILL51680x227240 (
);

FILL FILL_0__9884_ (
);

FILL FILL_0__9044_ (
);

AND2X2 _11735_ (
    .A(_1688_),
    .B(_1687_),
    .Y(_1653_[17])
);

AND2X2 _11315_ (
    .A(_1468_),
    .B(_1467_),
    .Y(_1455_[6])
);

FILL FILL331360x4940 (
);

FILL FILL_0__12811_ (
);

FILL FILL_1__16290_ (
);

FILL FILL209000x311220 (
);

FILL FILL_0__15283_ (
);

FILL FILL294120x266760 (
);

FILL FILL102600x256880 (
);

FILL FILL_1__8420_ (
);

FILL FILL83600x24700 (
);

FILL FILL350360x4940 (
);

FILL FILL_0__16488_ (
);

AND2X2 _16773_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_5707_)
);

AND2X2 _16353_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_5294_)
);

FILL FILL462080x74100 (
);

DFFSR _8695_ (
    .CLK(clk_bF$buf52),
    .D(_69_[13]),
    .Q(\datapath_1.regfile_1.regOut[2] [13]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL_1__10943_ (
);

BUFX2 BUFX2_insert370 (
    .A(_6321_),
    .Y(_6321__bF$buf0)
);

FILL FILL357200x306280 (
);

BUFX2 BUFX2_insert371 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf4 )
);

BUFX2 BUFX2_insert372 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf3 )
);

BUFX2 BUFX2_insert373 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf2 )
);

BUFX2 BUFX2_insert374 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf1 )
);

AND2X2 _17978_ (
    .A(_6236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_6895_)
);

BUFX2 BUFX2_insert375 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf0 )
);

AND2X2 _17558_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_6481_)
);

BUFX2 BUFX2_insert376 (
    .A(_6262_),
    .Y(_6262__bF$buf4)
);

OR2X2 _17138_ (
    .A(_6065_),
    .B(_6066_),
    .Y(_6067_)
);

BUFX2 BUFX2_insert377 (
    .A(_6262_),
    .Y(_6262__bF$buf3)
);

BUFX2 BUFX2_insert378 (
    .A(_6262_),
    .Y(_6262__bF$buf2)
);

AND2X2 _12693_ (
    .A(_2243_),
    .B(_2257_),
    .Y(_2258_)
);

BUFX2 BUFX2_insert379 (
    .A(_6262_),
    .Y(_6262__bF$buf1)
);

OR2X2 _12273_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[30] [25]),
    .Y(_1967_)
);

FILL FILL89680x167960 (
);

FILL FILL_0__18634_ (
);

FILL FILL291080x64220 (
);

FILL FILL_0__8735_ (
);

FILL FILL236360x59280 (
);

OR2X2 _13898_ (
    .A(\datapath_1.a [27]),
    .B(_3342__bF$buf2),
    .Y(_3332_)
);

AND2X2 _13478_ (
    .A(_3008_),
    .B(_3007_),
    .Y(\datapath_1.a3 [1])
);

AND2X2 _13058_ (
    .A(_2614_),
    .B(_2464_),
    .Y(_2615_)
);

FILL FILL47880x163020 (
);

FILL FILL_0__19419_ (
);

FILL FILL146680x266760 (
);

FILL FILL_0__14974_ (
);

FILL FILL_0__14134_ (
);

FILL FILL9120x138320 (
);

FILL FILL63840x19760 (
);

FILL FILL_1__11061_ (
);

FILL FILL_0__15759_ (
);

FILL FILL_0__15339_ (
);

OR2X2 _15624_ (
    .A(_4575_),
    .B(_4572_),
    .Y(_4576_)
);

OR2X2 _15204_ (
    .A(_4161_),
    .B(_4159_),
    .Y(_4162_)
);

FILL FILL186960x360620 (
);

FILL FILL_0__10474_ (
);

FILL FILL_0__10054_ (
);

AND2X2 _18096_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_7011_)
);

FILL FILL_0__16700_ (
);

FILL FILL400520x29640 (
);

FILL FILL9880x123500 (
);

FILL FILL_0__19172_ (
);

FILL FILL305520x113620 (
);

OR2X2 _16829_ (
    .A(_5761_),
    .B(_5760_),
    .Y(_5762_)
);

OR2X2 _16409_ (
    .A(_5333_),
    .B(_5348_),
    .Y(_5349_)
);

OR2X2 _11964_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_1801_)
);

FILL FILL_0__11259_ (
);

DFFSR _11544_ (
    .CLK(clk_bF$buf96),
    .D(_1521_[24]),
    .Q(\datapath_1.regfile_1.regOut[24] [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

OR2X2 _11124_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_1381_)
);

FILL FILL_0__17905_ (
);

FILL FILL_0__12200_ (
);

FILL FILL67640x19760 (
);

AND2X2 _12749_ (
    .A(_2311_),
    .B(_2313_),
    .Y(_2314_)
);

AND2X2 _12329_ (
    .A(_1984_),
    .B(_2047_),
    .Y(_1983_[0])
);

FILL FILL252320x355680 (
);

FILL FILL_0__13825_ (
);

FILL FILL_0__13405_ (
);

FILL FILL453720x108680 (
);

FILL FILL18240x83980 (
);

AND2X2 _16582_ (
    .A(_4135__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [21]),
    .Y(_5519_)
);

FILL FILL_0__16297_ (
);

AND2X2 _16162_ (
    .A(_4210__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_5106_)
);

FILL FILL_1__9014_ (
);

FILL FILL_1__10332_ (
);

FILL FILL275880x207480 (
);

OR2X2 _17787_ (
    .A(_6706_),
    .B(_6705_),
    .Y(_6707_)
);

FILL FILL352640x172900 (
);

AND2X2 _17367_ (
    .A(_6243_),
    .B(\datapath_1.PCJump_27_bF$buf0 ),
    .Y(_6293_)
);

FILL FILL_1__19450_ (
);

OR2X2 _12082_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_1916__bF$buf0),
    .Y(_1860_)
);

FILL FILL315400x4940 (
);

FILL FILL_0__18023_ (
);

OR2X2 _9289_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_464__bF$buf0),
    .Y(_438_)
);

FILL FILL484880x306280 (
);

OR2X2 _10815_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_1215_)
);

NAND2X1 _13287_ (
    .A(_2229_),
    .B(_2231_),
    .Y(_2830_)
);

FILL FILL122360x182780 (
);

FILL FILL_1__15790_ (
);

FILL FILL370120x9880 (
);

AND2X2 _19513_ (
    .A(_8377_),
    .B(_8376_),
    .Y(_8320_[28])
);

FILL FILL_0__9749_ (
);

FILL FILL278920x29640 (
);

FILL FILL462840x29640 (
);

FILL FILL_1__16155_ (
);

FILL FILL353400x4940 (
);

FILL FILL_0__15988_ (
);

AND2X2 _15853_ (
    .A(_4177__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_4802_)
);

OR2X2 _15433_ (
    .A(_4380_),
    .B(_4387_),
    .Y(_4388_)
);

FILL FILL246240x113620 (
);

INVX1 _15013_ (
    .A(\datapath_1.a3 [0]),
    .Y(_4002_)
);

FILL FILL_0__10283_ (
);

FILL FILL208240x0 (
);

FILL FILL45600x227240 (
);

FILL FILL432440x128440 (
);

FILL FILL368600x301340 (
);

FILL FILL176320x118560 (
);

FILL FILL349600x138320 (
);

FILL FILL_1__12495_ (
);

FILL FILL175560x44460 (
);

AND2X2 _16638_ (
    .A(_4210__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_5574_)
);

AND2X2 _16218_ (
    .A(_4142__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_5161_)
);

FILL FILL_0__11488_ (
);

OR2X2 _11773_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_1718__bF$buf4),
    .Y(_1714_)
);

FILL FILL_1__18301_ (
);

OR2X2 _11353_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .B(_1520__bF$buf0),
    .Y(_1494_)
);

FILL FILL_0__11068_ (
);

FILL FILL427880x247000 (
);

FILL FILL256120x0 (
);

OR2X2 _9921_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_759_)
);

OR2X2 _9501_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_539_)
);

FILL FILL119320x24700 (
);

FILL FILL394440x108680 (
);

FILL FILL303240x24700 (
);

NAND2X1 _12978_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(_2344_),
    .Y(_2539_)
);

AND2X2 _12558_ (
    .A(_2128_),
    .B(_2078_),
    .Y(_2079_)
);

OR2X2 _12138_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_1897_)
);

FILL FILL_0__18919_ (
);

FILL FILL_0__13634_ (
);

FILL FILL106400x247000 (
);

FILL FILL_0__13214_ (
);

FILL FILL386840x44460 (
);

OR2X2 _16391_ (
    .A(_5329_),
    .B(_5330_),
    .Y(_5331_)
);

FILL FILL179360x44460 (
);

FILL FILL206720x340860 (
);

FILL FILL_1__10141_ (
);

FILL FILL424840x143260 (
);

AND2X2 _14704_ (
    .A(_3855_),
    .B(_3854_),
    .Y(_3804_[25])
);

FILL FILL_0__14419_ (
);

FILL FILL199120x59280 (
);

BUFX2 BUFX2_insert750 (
    .A(_1520_),
    .Y(_1520__bF$buf2)
);

FILL FILL383040x59280 (
);

BUFX2 BUFX2_insert751 (
    .A(_1520_),
    .Y(_1520__bF$buf1)
);

BUFX2 BUFX2_insert752 (
    .A(_1520_),
    .Y(_1520__bF$buf0)
);

BUFX2 BUFX2_insert753 (
    .A(_6232_),
    .Y(_6232__bF$buf4)
);

BUFX2 BUFX2_insert754 (
    .A(_6232_),
    .Y(_6232__bF$buf3)
);

OR2X2 _17596_ (
    .A(_6517_),
    .B(_6518_),
    .Y(_6519_)
);

BUFX2 BUFX2_insert755 (
    .A(_6232_),
    .Y(_6232__bF$buf2)
);

FILL FILL488680x39520 (
);

BUFX2 BUFX2_insert756 (
    .A(_6232_),
    .Y(_6232__bF$buf1)
);

OR2X2 _17176_ (
    .A(_6103_),
    .B(_6096_),
    .Y(_6104_)
);

BUFX2 BUFX2_insert757 (
    .A(_6232_),
    .Y(_6232__bF$buf0)
);

BUFX2 BUFX2_insert758 (
    .A(_1652_),
    .Y(_1652__bF$buf4)
);

BUFX2 BUFX2_insert759 (
    .A(_1652_),
    .Y(_1652__bF$buf3)
);

FILL FILL324520x237120 (
);

FILL FILL_0__18672_ (
);

FILL FILL_0__18252_ (
);

FILL FILL223440x256880 (
);

DFFSR _9098_ (
    .CLK(clk_bF$buf0),
    .D(_267_[29]),
    .Q(\datapath_1.regfile_1.regOut[5] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

AND2X2 _15909_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_4857_)
);

FILL FILL347320x321100 (
);

FILL FILL_0__8773_ (
);

FILL FILL_0__10339_ (
);

DFFSR _10624_ (
    .CLK(clk_bF$buf39),
    .D(_1059_[7]),
    .Q(\datapath_1.regfile_1.regOut[17] [7]),
    .R(rst_bF$buf3),
    .S(vdd)
);

OR2X2 _10204_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .B(_926__bF$buf4),
    .Y(_908_)
);

FILL FILL240920x266760 (
);

FILL FILL310080x167960 (
);

OR2X2 _13096_ (
    .A(_2649_),
    .B(_2650_),
    .Y(_2651_)
);

FILL FILL_0__19457_ (
);

FILL FILL_0__19037_ (
);

OR2X2 _19322_ (
    .A(_8217_),
    .B(_8216_),
    .Y(_8218_)
);

FILL FILL172520x148200 (
);

FILL FILL_0__14592_ (
);

FILL FILL428640x251940 (
);

FILL FILL_0__9558_ (
);

FILL FILL_0__9138_ (
);

OR2X2 _11829_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_1731_)
);

DFFSR _11409_ (
    .CLK(clk_bF$buf3),
    .D(_1455_[18]),
    .Q(\datapath_1.regfile_1.regOut[23] [18]),
    .R(rst_bF$buf58),
    .S(vdd)
);

FILL FILL_0__12905_ (
);

FILL FILL_0__15377_ (
);

OR2X2 _15662_ (
    .A(_4612_),
    .B(_4613_),
    .Y(_4614_)
);

AND2X2 _15242_ (
    .A(_4166_),
    .B(_4144_),
    .Y(_4200_)
);

FILL FILL_0__10092_ (
);

OR2X2 _16867_ (
    .A(_5798_),
    .B(_5799_),
    .Y(_5800_)
);

FILL FILL348840x74100 (
);

AND2X2 _16447_ (
    .A(_4225__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_5386_)
);

AND2X2 _16027_ (
    .A(_4208__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_4973_)
);

FILL FILL_1__18950_ (
);

AND2X2 _11582_ (
    .A(_1606_),
    .B(_1605_),
    .Y(_1587_[9])
);

DFFSR _11162_ (
    .CLK(clk_bF$buf64),
    .D(_1323_[29]),
    .Q(\datapath_1.regfile_1.regOut[21] [29]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL_0__17943_ (
);

FILL FILL_0__17523_ (
);

FILL FILL_0__17103_ (
);

FILL FILL12920x207480 (
);

AND2X2 _8789_ (
    .A(_184_),
    .B(_183_),
    .Y(_135_[24])
);

FILL FILL115520x365560 (
);

DFFSR _9730_ (
    .CLK(clk_bF$buf0),
    .D(_597_[16]),
    .Q(\datapath_1.regfile_1.regOut[10] [16]),
    .R(rst_bF$buf64),
    .S(vdd)
);

OR2X2 _9310_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_464__bF$buf4),
    .Y(_452_)
);

INVX1 _12787_ (
    .A(\datapath_1.alu_1.ALUInB [29]),
    .Y(_2352_)
);

OR2X2 _12367_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .B(_2048__bF$buf3),
    .Y(_2010_)
);

FILL FILL_1__19315_ (
);

FILL FILL_1__14450_ (
);

FILL FILL348080x133380 (
);

FILL FILL_1__14030_ (
);

FILL FILL339720x202540 (
);

FILL FILL_0__13863_ (
);

FILL FILL_0__13023_ (
);

FILL FILL207480x34580 (
);

FILL FILL194560x14820 (
);

FILL FILL10640x59280 (
);

FILL FILL39520x212420 (
);

FILL FILL426360x113620 (
);

FILL FILL_1__9052_ (
);

FILL FILL_1__15655_ (
);

FILL FILL270560x103740 (
);

OR2X2 _14933_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [16]),
    .Y(_3968_)
);

FILL FILL_0__14648_ (
);

FILL FILL_0__14228_ (
);

OR2X2 _14513_ (
    .A(IRWrite_bF$buf3),
    .B(\aluControl_1.inst [5]),
    .Y(_3748_)
);

FILL FILL50920x375440 (
);

FILL FILL_0__18061_ (
);

FILL FILL_1__11995_ (
);

FILL FILL354920x286520 (
);

OR2X2 _15718_ (
    .A(_4667_),
    .B(_4668_),
    .Y(_4669_)
);

FILL FILL_0__10988_ (
);

AND2X2 _10853_ (
    .A(_1240_),
    .B(_1239_),
    .Y(_1191_[24])
);

AND2X2 _10433_ (
    .A(_1020_),
    .B(_1019_),
    .Y(_993_[13])
);

FILL FILL_0__10148_ (
);

AND2X2 _10013_ (
    .A(_800_),
    .B(_799_),
    .Y(_795_[2])
);

FILL FILL418000x143260 (
);

DFFSR _19551_ (
    .CLK(clk_bF$buf22),
    .D(_8320_[28]),
    .Q(\datapath_1.regfile_1.regOut[0] [28]),
    .R(rst_bF$buf7),
    .S(vdd)
);

FILL FILL_0__19266_ (
);

FILL FILL185440x187720 (
);

AND2X2 _19131_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_8030_)
);

FILL FILL_0__9787_ (
);

FILL FILL_0__9367_ (
);

OR2X2 _11638_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_1652__bF$buf2),
    .Y(_1644_)
);

OR2X2 _11218_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .B(_1454__bF$buf4),
    .Y(_1424_)
);

FILL FILL14440x311220 (
);

OR2X2 _15891_ (
    .A(_4838_),
    .B(_4837_),
    .Y(_4839_)
);

OR2X2 _15471_ (
    .A(_4422_),
    .B(_4425_),
    .Y(_4426_)
);

AND2X2 _15051_ (
    .A(_4039_),
    .B(_4037_),
    .Y(_4040_)
);

FILL FILL_1__8743_ (
);

FILL FILL_1__14506_ (
);

FILL FILL162640x212420 (
);

FILL FILL329840x291460 (
);

FILL FILL266000x24700 (
);

FILL FILL31160x227240 (
);

AND2X2 _16676_ (
    .A(_4195__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_5612_)
);

OR2X2 _16256_ (
    .A(_5197_),
    .B(_5196_),
    .Y(_5198_)
);

DFFSR _11391_ (
    .CLK(clk_bF$buf19),
    .D(_1455_[0]),
    .Q(\datapath_1.regfile_1.regOut[23] [0]),
    .R(rst_bF$buf19),
    .S(vdd)
);

FILL FILL_1__9948_ (
);

FILL FILL_0__17752_ (
);

OR2X2 _8598_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_77_)
);

FILL FILL134520x345800 (
);

FILL FILL315400x34580 (
);

FILL FILL160360x286520 (
);

FILL FILL205960x54340 (
);

INVX1 _12596_ (
    .A(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2161_)
);

DFFSR _12176_ (
    .CLK(clk_bF$buf57),
    .D(_1851_[11]),
    .Q(\datapath_1.regfile_1.regOut[29] [11]),
    .R(rst_bF$buf17),
    .S(vdd)
);

AND2X2 _18822_ (
    .A(_6287__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_7726_)
);

FILL FILL_0__18537_ (
);

FILL FILL_0__18117_ (
);

AND2X2 _18402_ (
    .A(_6300__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_7312_)
);

FILL FILL_0__13252_ (
);

FILL FILL_0__8638_ (
);

OR2X2 _10909_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(_1322__bF$buf3),
    .Y(_1258_)
);

FILL FILL_1__15884_ (
);

FILL FILL269800x345800 (
);

DFFSR _14742_ (
    .CLK(clk_bF$buf58),
    .D(_3804_[19]),
    .Q(\datapath_1.a [19]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__14457_ (
);

FILL FILL431680x4940 (
);

OR2X2 _14322_ (
    .A(\datapath_1.ALUResult [27]),
    .B(_3671__bF$buf2),
    .Y(_3661_)
);

FILL FILL171000x158080 (
);

FILL FILL319200x34580 (
);

FILL FILL_0__18290_ (
);

FILL FILL_1__11384_ (
);

AND2X2 _15947_ (
    .A(_4160__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_4894_)
);

OR2X2 _15527_ (
    .A(_4477_),
    .B(_4480_),
    .Y(_4481_)
);

AND2X2 _15107_ (
    .A(_4087_),
    .B(_4086_),
    .Y(_4088_)
);

FILL FILL284240x74100 (
);

FILL FILL_0__8391_ (
);

FILL FILL_0__10797_ (
);

OR2X2 _10662_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_1133_)
);

DFFSR _10242_ (
    .CLK(clk_bF$buf28),
    .D(_861_[12]),
    .Q(\datapath_1.regfile_1.regOut[14] [12]),
    .R(rst_bF$buf96),
    .S(vdd)
);

FILL FILL246240x19760 (
);

FILL FILL_0__16603_ (
);

FILL FILL_0__19495_ (
);

FILL FILL_0__19075_ (
);

AND2X2 _19360_ (
    .A(_8255_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd1 [30])
);

FILL FILL126160x266760 (
);

FILL FILL281200x113620 (
);

AND2X2 _8810_ (
    .A(_198_),
    .B(_197_),
    .Y(_135_[31])
);

FILL FILL448400x192660 (
);

FILL FILL_1__18815_ (
);

AND2X2 _11867_ (
    .A(_1756_),
    .B(_1755_),
    .Y(_1719_[18])
);

FILL FILL_0__9176_ (
);

AND2X2 _11447_ (
    .A(_1536_),
    .B(_1535_),
    .Y(_1521_[7])
);

DFFSR _11027_ (
    .CLK(clk_bF$buf26),
    .D(_1257_[23]),
    .Q(\datapath_1.regfile_1.regOut[20] [23]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL308560x177840 (
);

FILL FILL_0__12943_ (
);

FILL FILL_0__12523_ (
);

FILL FILL_0__12103_ (
);

OR2X2 _15280_ (
    .A(_4237_),
    .B(_4235_),
    .Y(_4238_)
);

FILL FILL44840x360620 (
);

FILL FILL_0__13728_ (
);

FILL FILL361760x266760 (
);

FILL FILL_0_BUFX2_insert1090 (
);

FILL FILL_0_BUFX2_insert1091 (
);

FILL FILL_0_BUFX2_insert1093 (
);

AND2X2 _16485_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_5424_)
);

OR2X2 _16065_ (
    .A(_5006_),
    .B(_5009_),
    .Y(_5010_)
);

FILL FILL_0_BUFX2_insert1095 (
);

FILL FILL_0_BUFX2_insert1097 (
);

FILL FILL_1__9757_ (
);

FILL FILL_0_BUFX2_insert1099 (
);

FILL FILL278920x276640 (
);

FILL FILL_0__17141_ (
);

FILL FILL106400x54340 (
);

FILL FILL505400x14820 (
);

FILL FILL20520x83980 (
);

FILL FILL_0__18766_ (
);

FILL FILL_0__18346_ (
);

AND2X2 _18631_ (
    .A(_6206__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_7538_)
);

AND2X2 _18211_ (
    .A(_6312__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_7124_)
);

FILL FILL342000x227240 (
);

FILL FILL_0__13481_ (
);

FILL FILL150480x163020 (
);

FILL FILL228000x251940 (
);

FILL FILL415720x49400 (
);

FILL FILL_0__8867_ (
);

FILL FILL_0__8447_ (
);

AND2X2 _10718_ (
    .A(_1170_),
    .B(_1169_),
    .Y(_1125_[22])
);

FILL FILL_1__12801_ (
);

FILL FILL_1__15273_ (
);

OR2X2 _19416_ (
    .A(_8309_),
    .B(_8310_),
    .Y(_8311_)
);

AND2X2 _14971_ (
    .A(_3993_),
    .B(_3992_),
    .Y(_3936_[28])
);

FILL FILL_0__14266_ (
);

AND2X2 _14551_ (
    .A(_3773_),
    .B(_3772_),
    .Y(_3738_[17])
);

AND2X2 _14131_ (
    .A(_3350__bF$buf2),
    .B(_2_[30]),
    .Y(_3532_)
);

FILL FILL475760x69160 (
);

FILL FILL_1__11193_ (
);

OR2X2 _15756_ (
    .A(_4705_),
    .B(_4704_),
    .Y(_4706_)
);

OR2X2 _15336_ (
    .A(_4292_),
    .B(_4285_),
    .Y(_4293_)
);

DFFSR _10891_ (
    .CLK(clk_bF$buf53),
    .D(_1191_[16]),
    .Q(\datapath_1.regfile_1.regOut[19] [16]),
    .R(rst_bF$buf111),
    .S(vdd)
);

OR2X2 _10471_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .B(_1058__bF$buf4),
    .Y(_1046_)
);

FILL FILL_0__10186_ (
);

OR2X2 _10051_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .B(_860__bF$buf3),
    .Y(_826_)
);

FILL FILL419520x49400 (
);

FILL FILL_0__16412_ (
);

FILL FILL_1__12398_ (
);

FILL FILL490960x207480 (
);

FILL FILL141360x54340 (
);

DFFSR _11676_ (
    .CLK(clk_bF$buf14),
    .D(_1587_[27]),
    .Q(\datapath_1.regfile_1.regOut[25] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

OR2X2 _11256_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_1449_)
);

FILL FILL_0__17617_ (
);

OR2X2 _17902_ (
    .A(_6819_),
    .B(_6818_),
    .Y(_6820_)
);

FILL FILL_0__12752_ (
);

FILL FILL_0__12332_ (
);

FILL FILL161120x69160 (
);

FILL FILL338200x163020 (
);

AND2X2 _9824_ (
    .A(_714_),
    .B(_713_),
    .Y(_663_[25])
);

AND2X2 _9404_ (
    .A(_494_),
    .B(_493_),
    .Y(_465_[14])
);

FILL FILL116280x330980 (
);

FILL FILL_1__14124_ (
);

OR2X2 _13822_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [2]),
    .Y(_3281_)
);

FILL FILL234840x321100 (
);

FILL FILL_0__13117_ (
);

OR2X2 _13402_ (
    .A(_2392_),
    .B(_2503_),
    .Y(_2938_)
);

OR2X2 _16294_ (
    .A(_5234_),
    .B(_5235_),
    .Y(_5236_)
);

FILL FILL82840x83980 (
);

FILL FILL_1__9146_ (
);

FILL FILL_0__17790_ (
);

FILL FILL_0__17370_ (
);

FILL FILL114760x177840 (
);

FILL FILL_1__15749_ (
);

FILL FILL_1__10464_ (
);

DFFSR _14607_ (
    .CLK(clk_bF$buf23),
    .D(_3738_[13]),
    .Q(\datapath_1.PCJump [15]),
    .R(rst_bF$buf33),
    .S(vdd)
);

OR2X2 _17499_ (
    .A(_6422_),
    .B(_6421_),
    .Y(_6423_)
);

OR2X2 _17079_ (
    .A(_6008_),
    .B(_6001_),
    .Y(_6009_)
);

FILL FILL_0__18995_ (
);

FILL FILL15960x261820 (
);

FILL FILL_0__18575_ (
);

OR2X2 _18860_ (
    .A(_7759_),
    .B(_7762_),
    .Y(_7763_)
);

AND2X2 _18440_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_7350_)
);

AND2X2 _18020_ (
    .A(_6264__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_6936_)
);

FILL FILL196080x207480 (
);

OR2X2 _10947_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_1283_)
);

OR2X2 _10527_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_1063_)
);

DFFSR _10107_ (
    .CLK(clk_bF$buf36),
    .D(_795_[6]),
    .Q(\datapath_1.regfile_1.regOut[13] [6]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL_0__11603_ (
);

FILL FILL490960x39520 (
);

OR2X2 _19225_ (
    .A(_8119_),
    .B(_8122_),
    .Y(_8123_)
);

OR2X2 _14780_ (
    .A(vdd),
    .B(_2_[8]),
    .Y(_3886_)
);

FILL FILL_0__14075_ (
);

DFFSR _14360_ (
    .CLK(clk_bF$buf20),
    .D(_3606_[24]),
    .Q(ALUOut[24]),
    .R(rst_bF$buf22),
    .S(vdd)
);

FILL FILL395200x360620 (
);

FILL FILL_0__12808_ (
);

AND2X2 _15985_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_4932_)
);

AND2X2 _15565_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_4518_)
);

INVX1 _15145_ (
    .A(_4111_),
    .Y(_4112_)
);

AND2X2 _10280_ (
    .A(_938_),
    .B(_937_),
    .Y(_927_[5])
);

FILL FILL_0__16641_ (
);

FILL FILL_0__16221_ (
);

FILL FILL266000x217360 (
);

OR2X2 _11485_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .B(_1586__bF$buf2),
    .Y(_1562_)
);

FILL FILL_1__18433_ (
);

OR2X2 _11065_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .B(_1388__bF$buf0),
    .Y(_1342_)
);

OR2X2 _17711_ (
    .A(_6630_),
    .B(_6631_),
    .Y(_6632_)
);

FILL FILL_0__17006_ (
);

FILL FILL_0__12981_ (
);

FILL FILL_0__12561_ (
);

FILL FILL13680x123500 (
);

OR2X2 _9633_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_607_)
);

DFFSR _9213_ (
    .CLK(clk_bF$buf17),
    .D(_333_[15]),
    .Q(\datapath_1.regfile_1.regOut[6] [15]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _18916_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_7818_)
);

FILL FILL503880x370500 (
);

FILL FILL_0__13766_ (
);

FILL FILL_0__13346_ (
);

OR2X2 _13631_ (
    .A(_3120_),
    .B(_3119_),
    .Y(_3121_)
);

OAI21X1 _13211_ (
    .A(_2755_),
    .B(_2501_),
    .C(_2758_),
    .Y(_2759_)
);

FILL FILL_1__15138_ (
);

FILL FILL_1__10273_ (
);

AND2X2 _14836_ (
    .A(_3923_),
    .B(_3922_),
    .Y(_3870_[26])
);

AND2X2 _14416_ (
    .A(_3703_),
    .B(_3702_),
    .Y(_3672_[15])
);

FILL FILL264480x276640 (
);

FILL FILL_0__15912_ (
);

FILL FILL_1__19391_ (
);

FILL FILL_0__18384_ (
);

FILL FILL_0__8485_ (
);

DFFSR _10756_ (
    .CLK(clk_bF$buf88),
    .D(_1125_[10]),
    .Q(\datapath_1.regfile_1.regOut[18] [10]),
    .R(rst_bF$buf95),
    .S(vdd)
);

OR2X2 _10336_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .B(_992__bF$buf3),
    .Y(_976_)
);

FILL FILL313120x355680 (
);

FILL FILL400520x360620 (
);

OR2X2 _19454_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [9]),
    .Y(_8338_)
);

OR2X2 _19034_ (
    .A(_7900_),
    .B(_7934_),
    .Y(_7935_)
);

OR2X2 _8904_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_241_)
);

FILL FILL327560x316160 (
);

FILL FILL414960x321100 (
);

FILL FILL_1__18909_ (
);

FILL FILL_1__13624_ (
);

FILL FILL_1_BUFX2_insert321 (
);

AND2X2 _12902_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2467_)
);

FILL FILL_0__12617_ (
);

FILL FILL_1_BUFX2_insert323 (
);

FILL FILL_1__16096_ (
);

FILL FILL_1_BUFX2_insert325 (
);

FILL FILL245480x222300 (
);

OR2X2 _15794_ (
    .A(_4742_),
    .B(_4743_),
    .Y(_4744_)
);

FILL FILL_0__15089_ (
);

AND2X2 _15374_ (
    .A(_4208__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_4330_)
);

FILL FILL_0__16870_ (
);

FILL FILL_1__14829_ (
);

FILL FILL385320x103740 (
);

FILL FILL408120x59280 (
);

FILL FILL376960x301340 (
);

OR2X2 _16999_ (
    .A(_5929_),
    .B(_5926_),
    .Y(_5930_)
);

AND2X2 _16579_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_5516_)
);

OR2X2 _16159_ (
    .A(_5101_),
    .B(_5102_),
    .Y(_5103_)
);

OR2X2 _11294_ (
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .Y(_1519_)
);

FILL FILL76760x311220 (
);

OR2X2 _17940_ (
    .A(_6856_),
    .B(_6855_),
    .Y(_6857_)
);

FILL FILL_0__17655_ (
);

FILL FILL_0__17235_ (
);

OR2X2 _17520_ (
    .A(_6440_),
    .B(_6443_),
    .Y(_6444_)
);

OR2X2 _17100_ (
    .A(_6028_),
    .B(_6027_),
    .Y(_6029_)
);

FILL FILL296400x266760 (
);

FILL FILL_0__12370_ (
);

FILL FILL66120x271700 (
);

FILL FILL480320x88920 (
);

FILL FILL167960x19760 (
);

DFFSR _9862_ (
    .CLK(clk_bF$buf86),
    .D(_663_[19]),
    .Q(\datapath_1.regfile_1.regOut[11] [19]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9442_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .B(_530__bF$buf2),
    .Y(_520_)
);

OR2X2 _9022_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .B(_332__bF$buf2),
    .Y(_300_)
);

AND2X2 _12499_ (
    .A(ALUSrcB[0]),
    .B(_2091_),
    .Y(IRWrite)
);

OR2X2 _12079_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .B(_1916__bF$buf0),
    .Y(_1858_)
);

FILL FILL_1__14582_ (
);

OR2X2 _18725_ (
    .A(_7626_),
    .B(_7629_),
    .Y(_7630_)
);

FILL FILL435480x345800 (
);

AND2X2 _18305_ (
    .A(_6250__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_7217_)
);

FILL FILL_0__13995_ (
);

FILL FILL179360x335920 (
);

AND2X2 _13860_ (
    .A(_3306_),
    .B(_3305_),
    .Y(\datapath_1.alu_1.ALUInA [14])
);

FILL FILL_0__13575_ (
);

INVX1 _13440_ (
    .A(_2973_),
    .Y(\datapath_1.ALUResult [0])
);

OAI21X1 _13020_ (
    .A(_2330_),
    .B(_2503_),
    .C(_2578_),
    .Y(_2579_)
);

FILL FILL114760x247000 (
);

FILL FILL237120x118560 (
);

FILL FILL_1__9184_ (
);

FILL FILL31920x281580 (
);

FILL FILL_1__10082_ (
);

OR2X2 _14645_ (
    .A(vdd),
    .B(\datapath_1.a [6]),
    .Y(_3816_)
);

OR2X2 _14225_ (
    .A(\datapath_1.Data [27]),
    .B(_3605__bF$buf3),
    .Y(_3595_)
);

FILL FILL345800x330980 (
);

FILL FILL110200x34580 (
);

FILL FILL_0__15721_ (
);

FILL FILL237880x103740 (
);

FILL FILL_0__18193_ (
);

FILL FILL218880x261820 (
);

FILL FILL_1__17933_ (
);

AND2X2 _10985_ (
    .A(_1308_),
    .B(_1307_),
    .Y(_1257_[25])
);

AND2X2 _10565_ (
    .A(_1088_),
    .B(_1087_),
    .Y(_1059_[14])
);

FILL FILL_1__17513_ (
);

AND2X2 _10145_ (
    .A(_868_),
    .B(_867_),
    .Y(_861_[3])
);

FILL FILL_0__16506_ (
);

FILL FILL_0__11221_ (
);

AND2X2 _19263_ (
    .A(_6323__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_8160_)
);

FILL FILL285760x326040 (
);

DFFSR _8713_ (
    .CLK(clk_bF$buf10),
    .D(_69_[31]),
    .Q(\datapath_1.regfile_1.regOut[2] [31]),
    .R(rst_bF$buf16),
    .S(vdd)
);

FILL FILL_0__9499_ (
);

FILL FILL_1__13013_ (
);

FILL FILL_0__12846_ (
);

OR2X2 _12711_ (
    .A(_2268_),
    .B(_2275_),
    .Y(_2276_)
);

FILL FILL_0__12006_ (
);

NOR2X1 _15183_ (
    .A(_4140_),
    .B(\datapath_1.PCJump_22_bF$buf0 ),
    .Y(_4141_)
);

FILL FILL63080x19760 (
);

OR2X2 _9918_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_757_)
);

FILL FILL_1__8875_ (
);

FILL FILL_1__14638_ (
);

FILL FILL66880x266760 (
);

AND2X2 _13916_ (
    .A(_3346_),
    .B(ALUSrcB[1]),
    .Y(_3347_)
);

OR2X2 _16388_ (
    .A(_5326_),
    .B(_5327_),
    .Y(_5328_)
);

FILL FILL_0__17884_ (
);

FILL FILL_0__17464_ (
);

FILL FILL_0__17044_ (
);

AND2X2 _9671_ (
    .A(_632_),
    .B(_631_),
    .Y(_597_[17])
);

AND2X2 _9251_ (
    .A(_412_),
    .B(_411_),
    .Y(_399_[6])
);

FILL FILL_1__19256_ (
);

FILL FILL_0__10912_ (
);

FILL FILL_1__14391_ (
);

AND2X2 _18954_ (
    .A(_6287__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_7856_)
);

AND2X2 _18534_ (
    .A(_6250__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_7442_)
);

AND2X2 _18114_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_7029_)
);

FILL FILL_0__13384_ (
);

FILL FILL364040x0 (
);

FILL FILL_0__9711_ (
);

OR2X2 _19319_ (
    .A(_8213_),
    .B(_8214_),
    .Y(_8215_)
);

FILL FILL354920x172900 (
);

DFFSR _14874_ (
    .CLK(clk_bF$buf98),
    .D(_3870_[22]),
    .Q(_2_[22]),
    .R(rst_bF$buf61),
    .S(vdd)
);

FILL FILL_0__14589_ (
);

FILL FILL_0__14169_ (
);

OR2X2 _14454_ (
    .A(memoryOutData[28]),
    .B(_3737__bF$buf0),
    .Y(_3729_)
);

AND2X2 _14034_ (
    .A(_3352__bF$buf1),
    .B(\datapath_1.PCJump [16]),
    .Y(_3449_)
);

FILL FILL459040x256880 (
);

FILL FILL_0__15530_ (
);

FILL FILL274360x29640 (
);

FILL FILL_0__15110_ (
);

FILL FILL180880x375440 (
);

FILL FILL390640x251940 (
);

FILL FILL210520x49400 (
);

OR2X2 _15659_ (
    .A(_4610_),
    .B(_4609_),
    .Y(_4611_)
);

AND2X2 _15239_ (
    .A(_4186_),
    .B(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_4197_)
);

OR2X2 _10794_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_1201_)
);

FILL FILL_0__10089_ (
);

DFFSR _10374_ (
    .CLK(clk_bF$buf112),
    .D(_927_[15]),
    .Q(\datapath_1.regfile_1.regOut[15] [15]),
    .R(rst_bF$buf113),
    .S(vdd)
);

FILL FILL_0__16735_ (
);

FILL FILL167960x4940 (
);

OR2X2 _16600_ (
    .A(_5529_),
    .B(_5536_),
    .Y(_5537_)
);

AND2X2 _19492_ (
    .A(_8363_),
    .B(_8362_),
    .Y(_8320_[21])
);

OR2X2 _19072_ (
    .A(_7971_),
    .B(_7970_),
    .Y(_7972_)
);

FILL FILL130720x64220 (
);

DFFSR _8942_ (
    .CLK(clk_bF$buf111),
    .D(_201_[2]),
    .Q(\datapath_1.regfile_1.regOut[4] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

AND2X2 _8522_ (
    .A(_46_),
    .B(_45_),
    .Y(_3_[21])
);

FILL FILL359480x335920 (
);

FILL FILL500080x108680 (
);

AND2X2 _11999_ (
    .A(_1824_),
    .B(_1823_),
    .Y(_1785_[19])
);

AND2X2 _11579_ (
    .A(_1604_),
    .B(_1603_),
    .Y(_1587_[8])
);

DFFSR _11159_ (
    .CLK(clk_bF$buf54),
    .D(_1323_[26]),
    .Q(\datapath_1.regfile_1.regOut[21] [26]),
    .R(rst_bF$buf24),
    .S(vdd)
);

FILL FILL_1__13662_ (
);

FILL FILL_1__13242_ (
);

NOR2X1 _17805_ (
    .A(_6310__bF$buf0),
    .B(_6723_),
    .Y(_6724_)
);

FILL FILL_1_BUFX2_insert701 (
);

FILL FILL278160x29640 (
);

INVX1 _12940_ (
    .A(_2503_),
    .Y(_2504_)
);

FILL FILL_1_BUFX2_insert703 (
);

FILL FILL_0__12235_ (
);

INVX1 _12520_ (
    .A(\control_1.op [2]),
    .Y(_2110_)
);

OR2X2 _12100_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .B(_1916__bF$buf1),
    .Y(_1872_)
);

FILL FILL_1_BUFX2_insert705 (
);

FILL FILL373920x158080 (
);

FILL FILL436240x93860 (
);

DFFSR _9727_ (
    .CLK(clk_bF$buf13),
    .D(_597_[13]),
    .Q(\datapath_1.regfile_1.regOut[10] [13]),
    .R(rst_bF$buf90),
    .S(vdd)
);

OR2X2 _9307_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .B(_464__bF$buf0),
    .Y(_450_)
);

FILL FILL178600x118560 (
);

FILL FILL91200x34580 (
);

AND2X2 _13725_ (
    .A(_3084__bF$buf0),
    .B(\datapath_1.PCJump [19]),
    .Y(_3201_)
);

AND2X2 _13305_ (
    .A(_2846_),
    .B(_2837_),
    .Y(_2847_)
);

FILL FILL256880x227240 (
);

AND2X2 _16197_ (
    .A(_4151__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_5140_)
);

FILL FILL_0__14801_ (
);

FILL FILL_1__9889_ (
);

FILL FILL_0__17693_ (
);

FILL FILL282720x360620 (
);

FILL FILL279680x311220 (
);

FILL FILL396720x108680 (
);

DFFSR _9480_ (
    .CLK(clk_bF$buf96),
    .D(_465_[24]),
    .Q(\datapath_1.regfile_1.regOut[8] [24]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9060_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_325_)
);

FILL FILL_1__19485_ (
);

FILL FILL455240x286520 (
);

FILL FILL_0__10301_ (
);

OR2X2 _18763_ (
    .A(_7664_),
    .B(_7667_),
    .Y(_7668_)
);

FILL FILL_0__18478_ (
);

AND2X2 _18343_ (
    .A(_6262__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_7254_)
);

FILL FILL_0__18058_ (
);

FILL FILL_0__13193_ (
);

FILL FILL178600x14820 (
);

FILL FILL_0__8999_ (
);

FILL FILL_0__9940_ (
);

FILL FILL476520x83980 (
);

FILL FILL_0__11506_ (
);

FILL FILL340480x74100 (
);

FILL FILL272840x49400 (
);

DFFSR _19548_ (
    .CLK(clk_bF$buf69),
    .D(_8320_[25]),
    .Q(\datapath_1.regfile_1.regOut[0] [25]),
    .R(rst_bF$buf76),
    .S(vdd)
);

OR2X2 _19128_ (
    .A(_8019_),
    .B(_8026_),
    .Y(_8027_)
);

AND2X2 _14683_ (
    .A(_3841_),
    .B(_3840_),
    .Y(_3804_[18])
);

FILL FILL_0__14398_ (
);

AND2X2 _14263_ (
    .A(_3621_),
    .B(_3620_),
    .Y(_3606_[7])
);

FILL FILL326800x237120 (
);

FILL FILL225720x256880 (
);

FILL FILL240160x128440 (
);

FILL FILL413440x148200 (
);

FILL FILL349600x321100 (
);

OR2X2 _15888_ (
    .A(_4832_),
    .B(_4835_),
    .Y(_4836_)
);

AND2X2 _15468_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_4423_)
);

NAND3X1 _15048_ (
    .A(_4013_),
    .B(_4017_),
    .C(_4012_),
    .Y(_4037_)
);

FILL FILL_1__17551_ (
);

OR2X2 _10183_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .B(_926__bF$buf0),
    .Y(_894_)
);

FILL FILL_0__16124_ (
);

FILL FILL88920x133380 (
);

OR2X2 _8751_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_159_)
);

OR2X2 _11388_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_1517_)
);

FILL FILL_1__13891_ (
);

FILL FILL_0__17749_ (
);

AND2X2 _17614_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_6536_)
);

FILL FILL_0__17329_ (
);

FILL FILL_0__12884_ (
);

FILL FILL_0__12464_ (
);

FILL FILL466640x330980 (
);

AND2X2 _9956_ (
    .A(_782_),
    .B(_781_),
    .Y(_729_[26])
);

AND2X2 _9536_ (
    .A(_562_),
    .B(_561_),
    .Y(_531_[15])
);

AND2X2 _9116_ (
    .A(_342_),
    .B(_341_),
    .Y(_333_[4])
);

OR2X2 _18819_ (
    .A(_7722_),
    .B(_7721_),
    .Y(_7723_)
);

FILL FILL_0_BUFX2_insert360 (
);

FILL FILL_0_BUFX2_insert362 (
);

AND2X2 _13954_ (
    .A(_3347__bF$buf1),
    .B(\aluControl_1.inst [5]),
    .Y(_3380_)
);

FILL FILL_0_BUFX2_insert364 (
);

FILL FILL_0__13669_ (
);

FILL FILL_0__13249_ (
);

FILL FILL_0_BUFX2_insert365 (
);

OR2X2 _13534_ (
    .A(IorD_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [15]),
    .Y(_3044_)
);

AND2X2 _13114_ (
    .A(_2666_),
    .B(_2294_),
    .Y(_2667_)
);

FILL FILL_0_BUFX2_insert366 (
);

FILL FILL267520x0 (
);

FILL FILL_0_BUFX2_insert367 (
);

FILL FILL_0_BUFX2_insert368 (
);

FILL FILL117800x365560 (
);

FILL FILL_1__9278_ (
);

FILL FILL_0__17082_ (
);

DFFSR _14739_ (
    .CLK(clk_bF$buf15),
    .D(_3804_[16]),
    .Q(\datapath_1.a [16]),
    .R(rst_bF$buf91),
    .S(vdd)
);

OR2X2 _14319_ (
    .A(\datapath_1.ALUResult [26]),
    .B(_3671__bF$buf1),
    .Y(_3659_)
);

FILL FILL_1__16402_ (
);

FILL FILL_0__10950_ (
);

AND2X2 _18992_ (
    .A(_6259__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_7893_)
);

AND2X2 _18572_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_7480_)
);

OR2X2 _18152_ (
    .A(_7062_),
    .B(_7065_),
    .Y(_7066_)
);

FILL FILL253080x4940 (
);

FILL FILL428640x113620 (
);

FILL FILL158080x98800 (
);

OR2X2 _10659_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_1131_)
);

DFFSR _10239_ (
    .CLK(clk_bF$buf89),
    .D(_861_[9]),
    .Q(\datapath_1.regfile_1.regOut[14] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

FILL FILL_1__12742_ (
);

FILL FILL409640x271700 (
);

FILL FILL_0__11735_ (
);

FILL FILL35720x365560 (
);

AND2X2 _11600_ (
    .A(_1618_),
    .B(_1617_),
    .Y(_1587_[15])
);

FILL FILL_0__11315_ (
);

OR2X2 _19357_ (
    .A(_8252_),
    .B(_8237_),
    .Y(_8253_)
);

DFFSR _14492_ (
    .CLK(clk_bF$buf42),
    .D(_3672_[27]),
    .Q(\datapath_1.Data [27]),
    .R(rst_bF$buf100),
    .S(vdd)
);

AND2X2 _14072_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3481_)
);

FILL FILL272080x330980 (
);

AND2X2 _8807_ (
    .A(_196_),
    .B(_195_),
    .Y(_135_[30])
);

FILL FILL272080x4940 (
);

FILL FILL_1__13107_ (
);

FILL FILL426360x187720 (
);

OR2X2 _12805_ (
    .A(_2167_),
    .B(_2369_),
    .Y(_2370_)
);

FILL FILL369360x98800 (
);

AND2X2 _15697_ (
    .A(_4214__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_4648_)
);

AND2X2 _15277_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_4235_)
);

FILL FILL291080x4940 (
);

FILL FILL443840x197600 (
);

FILL FILL_0__16773_ (
);

FILL FILL_0__16353_ (
);

OR2X2 _8980_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_332__bF$buf3),
    .Y(_272_)
);

DFFSR _8560_ (
    .CLK(clk_bF$buf48),
    .D(_3_[7]),
    .Q(\datapath_1.regfile_1.regOut[1] [7]),
    .R(rst_bF$buf14),
    .S(vdd)
);

OR2X2 _11197_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .B(_1454__bF$buf4),
    .Y(_1410_)
);

FILL FILL_0__17978_ (
);

FILL FILL16720x311220 (
);

FILL FILL_0__17558_ (
);

AND2X2 _17843_ (
    .A(_6264__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_6762_)
);

OR2X2 _17423_ (
    .A(_6347_),
    .B(_6346_),
    .Y(_6348_)
);

OR2X2 _17003_ (
    .A(_5932_),
    .B(_5933_),
    .Y(_5934_)
);

FILL FILL_0__12693_ (
);

OR2X2 _9765_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_675_)
);

DFFSR _9345_ (
    .CLK(clk_bF$buf103),
    .D(_399_[18]),
    .Q(\datapath_1.regfile_1.regOut[7] [18]),
    .R(rst_bF$buf0),
    .S(vdd)
);

FILL FILL346560x163020 (
);

FILL FILL_1__14065_ (
);

AND2X2 _18628_ (
    .A(_6321__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_7535_)
);

AND2X2 _18208_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_7121_)
);

FILL FILL33440x227240 (
);

FILL FILL_0__13898_ (
);

FILL FILL119320x335920 (
);

FILL FILL418000x19760 (
);

AND2X2 _13763_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3234_)
);

FILL FILL_0__13058_ (
);

OAI21X1 _13343_ (
    .A(_2500_),
    .B(_2871_),
    .C(_2383_),
    .Y(_2883_)
);

FILL FILL382280x242060 (
);

AND2X2 _14968_ (
    .A(_3991_),
    .B(_3990_),
    .Y(_3936_[27])
);

FILL FILL162640x286520 (
);

AND2X2 _14548_ (
    .A(_3771_),
    .B(_3770_),
    .Y(_3738_[16])
);

AND2X2 _14128_ (
    .A(_3344__bF$buf1),
    .B(gnd),
    .Y(_3529_)
);

FILL FILL_1__16631_ (
);

FILL FILL_0__15624_ (
);

FILL FILL_0__15204_ (
);

FILL FILL382280x108680 (
);

FILL FILL_0__18096_ (
);

OR2X2 _18381_ (
    .A(_7284_),
    .B(_7291_),
    .Y(_7292_)
);

FILL FILL37240x335920 (
);

DFFSR _10888_ (
    .CLK(clk_bF$buf34),
    .D(_1191_[13]),
    .Q(\datapath_1.regfile_1.regOut[19] [13]),
    .R(rst_bF$buf51),
    .S(vdd)
);

OR2X2 _10468_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .B(_1058__bF$buf3),
    .Y(_1044_)
);

OR2X2 _10048_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .B(_860__bF$buf0),
    .Y(_824_)
);

FILL FILL_0__16829_ (
);

FILL FILL_0__11124_ (
);

AND2X2 _19166_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_8064_)
);

OR2X2 _8616_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_89_)
);

FILL FILL80560x286520 (
);

FILL FILL459800x69160 (
);

FILL FILL_1__13756_ (
);

FILL FILL384560x197600 (
);

FILL FILL_0__12749_ (
);

AND2X2 _12614_ (
    .A(_2178_),
    .B(\datapath_1.alu_1.ALUInB [0]),
    .Y(_2179_)
);

FILL FILL269040x19760 (
);

FILL FILL211280x256880 (
);

NAND3X1 _15086_ (
    .A(_4020_),
    .B(_4002_),
    .C(_4017_),
    .Y(_4071_)
);

FILL FILL_1__8778_ (
);

FILL FILL12160x247000 (
);

FILL FILL128440x266760 (
);

FILL FILL_0__16582_ (
);

FILL FILL_0__16162_ (
);

FILL FILL215840x271700 (
);

OR2X2 _13819_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [1]),
    .Y(_3279_)
);

FILL FILL475000x202540 (
);

FILL FILL_1__18374_ (
);

FILL FILL79800x29640 (
);

AND2X2 _17652_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [4]),
    .Y(_6574_)
);

OR2X2 _17232_ (
    .A(_6155_),
    .B(_6158_),
    .Y(_6159_)
);

FILL FILL_0__12082_ (
);

FILL FILL256120x4940 (
);

FILL FILL297160x301340 (
);

FILL FILL433960x261820 (
);

DFFSR _9994_ (
    .CLK(clk_bF$buf72),
    .D(_729_[22]),
    .Q(\datapath_1.regfile_1.regOut[12] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

OR2X2 _9574_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_596__bF$buf2),
    .Y(_588_)
);

OR2X2 _9154_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .B(_398__bF$buf4),
    .Y(_368_)
);

FILL FILL458280x79040 (
);

FILL FILL_0__10815_ (
);

AND2X2 _18857_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_7760_)
);

FILL FILL_0_BUFX2_insert741 (
);

OR2X2 _18437_ (
    .A(_7346_),
    .B(_7345_),
    .Y(_7347_)
);

AND2X2 _18017_ (
    .A(_6259__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_6933_)
);

FILL FILL_0_BUFX2_insert743 (
);

AND2X2 _13992_ (
    .A(_3352__bF$buf0),
    .B(\datapath_1.PCJump [10]),
    .Y(_3413_)
);

FILL FILL_0_BUFX2_insert744 (
);

FILL FILL_0__13287_ (
);

FILL FILL_0_BUFX2_insert745 (
);

AND2X2 _13572_ (
    .A(_3069_),
    .B(_3068_),
    .Y(_1_[27])
);

NOR2X1 _13152_ (
    .A(_2503_),
    .B(_2282_),
    .Y(_2703_)
);

FILL FILL_0_BUFX2_insert746 (
);

FILL FILL_0_BUFX2_insert747 (
);

FILL FILL_0_BUFX2_insert748 (
);

FILL FILL_0__19513_ (
);

FILL FILL_1__12607_ (
);

FILL FILL_1__15079_ (
);

FILL FILL357960x93860 (
);

OR2X2 _14777_ (
    .A(vdd),
    .B(_2_[7]),
    .Y(_3884_)
);

DFFSR _14357_ (
    .CLK(clk_bF$buf41),
    .D(_3606_[21]),
    .Q(ALUOut[21]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL_1__16020_ (
);

FILL FILL_0__15853_ (
);

FILL FILL78280x39520 (
);

FILL FILL240160x39520 (
);

FILL FILL120840x375440 (
);

AND2X2 _18190_ (
    .A(_7103_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd1 [12])
);

AND2X2 _10697_ (
    .A(_1156_),
    .B(_1155_),
    .Y(_1125_[15])
);

AND2X2 _10277_ (
    .A(_936_),
    .B(_935_),
    .Y(_927_[4])
);

FILL FILL_1__12780_ (
);

FILL FILL_0__16638_ (
);

AND2X2 _16923_ (
    .A(_4208__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_5855_)
);

OR2X2 _16503_ (
    .A(_5441_),
    .B(_5434_),
    .Y(_5442_)
);

FILL FILL_0__16218_ (
);

FILL FILL505400x88920 (
);

FILL FILL_0__11353_ (
);

AND2X2 _19395_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_8290_)
);

OR2X2 _8845_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(_266__bF$buf1),
    .Y(_202_)
);

BUFX2 _8425_ (
    .A(_2_[1]),
    .Y(memoryWriteData[1])
);

OR2X2 _17708_ (
    .A(_6628_),
    .B(_6625_),
    .Y(_6629_)
);

FILL FILL_0__12978_ (
);

OR2X2 _12843_ (
    .A(_2406_),
    .B(_2407_),
    .Y(_2408_)
);

FILL FILL_0__12558_ (
);

FILL FILL_0__12138_ (
);

DFFSR _12423_ (
    .CLK(clk_bF$buf105),
    .D(_1983_[0]),
    .Q(\datapath_1.regfile_1.regOut[31] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

OR2X2 _12003_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[28] [21]),
    .Y(_1827_)
);

FILL FILL342760x286520 (
);

FILL FILL_1__8587_ (
);

FILL FILL371640x54340 (
);

FILL FILL19000x242060 (
);

OR2X2 _13628_ (
    .A(_3116_),
    .B(_3117_),
    .Y(_3118_)
);

NAND2X1 _13208_ (
    .A(_2755_),
    .B(_2548_),
    .Y(_2756_)
);

FILL FILL250040x133380 (
);

FILL FILL_0__14704_ (
);

OR2X2 _17881_ (
    .A(_6798_),
    .B(_6790_),
    .Y(_6799_)
);

FILL FILL_0__17596_ (
);

AND2X2 _17461_ (
    .A(_6232__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_6386_)
);

FILL FILL_0__17176_ (
);

AND2X2 _17041_ (
    .A(_4203__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_5971_)
);

FILL FILL_1__16916_ (
);

AND2X2 _9383_ (
    .A(_480_),
    .B(_479_),
    .Y(_465_[7])
);

FILL FILL_0__10204_ (
);

OR2X2 _18666_ (
    .A(_7567_),
    .B(_7571_),
    .Y(_7572_)
);

OR2X2 _18246_ (
    .A(_7157_),
    .B(_7158_),
    .Y(_7159_)
);

INVX1 _13381_ (
    .A(_2918_),
    .Y(\datapath_1.ALUResult [4])
);

FILL FILL_0__19322_ (
);

FILL FILL277400x9880 (
);

FILL FILL_0__9423_ (
);

FILL FILL_0__11829_ (
);

FILL FILL_0__9003_ (
);

FILL FILL463600x113620 (
);

OR2X2 _14586_ (
    .A(memoryOutData[29]),
    .B(_3803__bF$buf3),
    .Y(_3797_)
);

FILL FILL6080x93860 (
);

AND2X2 _14166_ (
    .A(_3555_),
    .B(_3554_),
    .Y(\datapath_1.mux_wd3.dout [7])
);

FILL FILL367840x306280 (
);

FILL FILL_0__15242_ (
);

FILL FILL_1_BUFX2_insert296 (
);

FILL FILL_1_BUFX2_insert298 (
);

FILL FILL480320x350740 (
);

OR2X2 _10086_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_849_)
);

FILL FILL_0__16867_ (
);

FILL FILL34960x177840 (
);

OR2X2 _16732_ (
    .A(_5666_),
    .B(_5665_),
    .Y(_5667_)
);

FILL FILL_0__16447_ (
);

FILL FILL_0__16027_ (
);

OR2X2 _16312_ (
    .A(_5238_),
    .B(_5253_),
    .Y(_5254_)
);

FILL FILL133000x217360 (
);

FILL FILL205960x158080 (
);

FILL FILL494760x311220 (
);

AND2X2 _8654_ (
    .A(_114_),
    .B(_113_),
    .Y(_69_[22])
);

FILL FILL231800x291460 (
);

FILL FILL_1__18239_ (
);

OR2X2 _17937_ (
    .A(_6850_),
    .B(_6853_),
    .Y(_6854_)
);

AND2X2 _17517_ (
    .A(_6211__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_6441_)
);

FILL FILL_0__12787_ (
);

FILL FILL_0__12367_ (
);

OR2X2 _12652_ (
    .A(_2213_),
    .B(_2216_),
    .Y(_2217_)
);

OR2X2 _12232_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .B(_1982__bF$buf4),
    .Y(_1940_)
);

DFFSR _9859_ (
    .CLK(clk_bF$buf88),
    .D(_663_[16]),
    .Q(\datapath_1.regfile_1.regOut[11] [16]),
    .R(rst_bF$buf95),
    .S(vdd)
);

OR2X2 _9439_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_530__bF$buf4),
    .Y(_518_)
);

OR2X2 _9019_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_332__bF$buf3),
    .Y(_298_)
);

FILL FILL_1__8396_ (
);

FILL FILL107920x69160 (
);

AND2X2 _13857_ (
    .A(_3304_),
    .B(_3303_),
    .Y(\datapath_1.alu_1.ALUInA [13])
);

AND2X2 _13437_ (
    .A(_2969_),
    .B(_2970_),
    .Y(_2971_)
);

NOR2X1 _13017_ (
    .A(_2501_),
    .B(_2329_),
    .Y(_2576_)
);

FILL FILL_1__15520_ (
);

FILL FILL_1__15100_ (
);

FILL FILL_0__14933_ (
);

FILL FILL_0__14513_ (
);

OR2X2 _17690_ (
    .A(_6609_),
    .B(_6610_),
    .Y(_6611_)
);

OR2X2 _17270_ (
    .A(_6193_),
    .B(_6196_),
    .Y(_6197_)
);

OR2X2 _9192_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_393_)
);

FILL FILL_0__15718_ (
);

FILL FILL353400x296400 (
);

FILL FILL_0__10433_ (
);

FILL FILL_0__10013_ (
);

AND2X2 _18895_ (
    .A(_6300__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_7798_)
);

AND2X2 _18475_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_7384_)
);

OR2X2 _18055_ (
    .A(_6967_),
    .B(_6970_),
    .Y(_6971_)
);

NAND2X1 _13190_ (
    .A(_2416_),
    .B(_2504_),
    .Y(_2739_)
);

FILL FILL_0__19131_ (
);

FILL FILL_0__11638_ (
);

FILL FILL_0__9232_ (
);

DFFSR _11923_ (
    .CLK(clk_bF$buf11),
    .D(_1719_[16]),
    .Q(\datapath_1.regfile_1.regOut[27] [16]),
    .R(rst_bF$buf111),
    .S(vdd)
);

OR2X2 _11503_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .B(_1586__bF$buf4),
    .Y(_1574_)
);

AND2X2 _14395_ (
    .A(_3689_),
    .B(_3688_),
    .Y(_3672_[8])
);

FILL FILL_0__15891_ (
);

FILL FILL_0__15471_ (
);

FILL FILL_0__15051_ (
);

FILL FILL407360x44460 (
);

NAND2X1 _12708_ (
    .A(_2271_),
    .B(_2272_),
    .Y(_2273_)
);

FILL FILL_0__16676_ (
);

OR2X2 _16961_ (
    .A(_5888_),
    .B(_5891_),
    .Y(_5892_)
);

AND2X2 _16541_ (
    .A(_4228__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_5479_)
);

OR2X2 _16121_ (
    .A(_5065_),
    .B(_5034_),
    .Y(_5066_)
);

FILL FILL329840x316160 (
);

OR2X2 _8883_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_227_)
);

OR2X2 _8463_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_7_)
);

FILL FILL_1__18888_ (
);

FILL FILL_1__18468_ (
);

FILL FILL_1__13183_ (
);

INVX1 _17746_ (
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_6666_)
);

OR2X2 _17326_ (
    .A(_6248_),
    .B(_6251_),
    .Y(_6252_)
);

AND2X2 _12881_ (
    .A(_2445_),
    .B(_2416_),
    .Y(_2446_)
);

AND2X2 _12461_ (
    .A(_2054_),
    .B(ALUOp[1]),
    .Y(_2055_)
);

DFFSR _12041_ (
    .CLK(clk_bF$buf104),
    .D(_1785_[5]),
    .Q(\datapath_1.regfile_1.regOut[28] [5]),
    .R(rst_bF$buf25),
    .S(vdd)
);

FILL FILL38760x217360 (
);

FILL FILL_0__18402_ (
);

AND2X2 _9668_ (
    .A(_630_),
    .B(_629_),
    .Y(_597_[16])
);

FILL FILL241680x375440 (
);

AND2X2 _9248_ (
    .A(_410_),
    .B(_409_),
    .Y(_399_[5])
);

FILL FILL387600x103740 (
);

FILL FILL_0__8503_ (
);

OR2X2 _13666_ (
    .A(_3150_),
    .B(_3149_),
    .Y(_3151_)
);

OR2X2 _13246_ (
    .A(_2220_),
    .B(_2210_),
    .Y(_2791_)
);

FILL FILL381520x256880 (
);

FILL FILL_1_BUFX2_insert1056 (
);

FILL FILL_1_BUFX2_insert1058 (
);

FILL FILL245480x296400 (
);

FILL FILL_0__14322_ (
);

FILL FILL_0__9708_ (
);

FILL FILL237120x0 (
);

FILL FILL304000x44460 (
);

FILL FILL_0__15947_ (
);

OR2X2 _15812_ (
    .A(_4760_),
    .B(_4759_),
    .Y(_4761_)
);

FILL FILL_0__15107_ (
);

OR2X2 _18284_ (
    .A(_7195_),
    .B(_7187_),
    .Y(_7196_)
);

FILL FILL214320x79040 (
);

FILL FILL294880x34580 (
);

FILL FILL239400x118560 (
);

FILL FILL_0__19360_ (
);

FILL FILL_1__17319_ (
);

FILL FILL_1__12874_ (
);

FILL FILL_1__12034_ (
);

FILL FILL_0__9881_ (
);

FILL FILL_0__11867_ (
);

FILL FILL152760x326040 (
);

FILL FILL_0__11447_ (
);

AND2X2 _11732_ (
    .A(_1686_),
    .B(_1685_),
    .Y(_1653_[16])
);

AND2X2 _11312_ (
    .A(_1466_),
    .B(_1465_),
    .Y(_1455_[5])
);

AND2X2 _19489_ (
    .A(_8361_),
    .B(_8360_),
    .Y(_8320_[20])
);

OR2X2 _19069_ (
    .A(_7967_),
    .B(_7968_),
    .Y(_7969_)
);

FILL FILL142120x286520 (
);

FILL FILL238640x14820 (
);

AND2X2 _8939_ (
    .A(_264_),
    .B(_263_),
    .Y(_201_[31])
);

AND2X2 _8519_ (
    .A(_44_),
    .B(_43_),
    .Y(_3_[20])
);

FILL FILL_0__15280_ (
);

FILL FILL474240x158080 (
);

FILL FILL332880x49400 (
);

NAND3X1 _12937_ (
    .A(_2386_),
    .B(_2500_),
    .C(ALUControl[0]),
    .Y(_2501_)
);

AND2X2 _12517_ (
    .A(ALUSrcB[0]),
    .B(\control_1.reg_state.dout [0]),
    .Y(_2108_)
);

FILL FILL366320x123500 (
);

FILL FILL_1_BUFX2_insert676 (
);

FILL FILL_1_BUFX2_insert678 (
);

FILL FILL334400x335920 (
);

FILL FILL34960x247000 (
);

FILL FILL218120x79040 (
);

FILL FILL_1__17492_ (
);

FILL FILL_1__17072_ (
);

AND2X2 _16770_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_5704_)
);

FILL FILL_0__16065_ (
);

AND2X2 _16350_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_5291_)
);

FILL FILL215840x88920 (
);

DFFSR _8692_ (
    .CLK(clk_bF$buf30),
    .D(_69_[10]),
    .Q(\datapath_1.regfile_1.regOut[2] [10]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL100320x148200 (
);

FILL FILL60040x286520 (
);

FILL FILL383040x360620 (
);

FILL FILL_1__10520_ (
);

FILL FILL497040x108680 (
);

BUFX2 BUFX2_insert340 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf1 )
);

BUFX2 BUFX2_insert341 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf0 )
);

BUFX2 BUFX2_insert342 (
    .A(_4234_),
    .Y(_4234__bF$buf4)
);

BUFX2 BUFX2_insert343 (
    .A(_4234_),
    .Y(_4234__bF$buf3)
);

BUFX2 BUFX2_insert344 (
    .A(_4234_),
    .Y(_4234__bF$buf2)
);

OR2X2 _17975_ (
    .A(_6891_),
    .B(_6884_),
    .Y(_6892_)
);

OR2X2 _17555_ (
    .A(_6470_),
    .B(_6477_),
    .Y(_6478_)
);

BUFX2 BUFX2_insert345 (
    .A(_4234_),
    .Y(_4234__bF$buf1)
);

BUFX2 BUFX2_insert346 (
    .A(_4234_),
    .Y(_4234__bF$buf0)
);

OR2X2 _17135_ (
    .A(_6063_),
    .B(_6060_),
    .Y(_6064_)
);

BUFX2 BUFX2_insert347 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf3 )
);

BUFX2 BUFX2_insert348 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf2 )
);

OR2X2 _12690_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(_2254_),
    .Y(_2255_)
);

BUFX2 BUFX2_insert349 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf1 )
);

OR2X2 _12270_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_1965_)
);

FILL FILL_0__18631_ (
);

FILL FILL_0__18211_ (
);

OR2X2 _9897_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_743_)
);

FILL FILL31920x143260 (
);

DFFSR _9477_ (
    .CLK(clk_bF$buf21),
    .D(_465_[21]),
    .Q(\datapath_1.regfile_1.regOut[8] [21]),
    .R(rst_bF$buf4),
    .S(vdd)
);

OR2X2 _9057_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_323_)
);

FILL FILL_1__11725_ (
);

FILL FILL495520x276640 (
);

FILL FILL_0__10718_ (
);

FILL FILL423320x316160 (
);

FILL FILL_1__14197_ (
);

FILL FILL254600x311220 (
);

OR2X2 _13895_ (
    .A(\datapath_1.a [26]),
    .B(_3342__bF$buf0),
    .Y(_3330_)
);

AND2X2 _13475_ (
    .A(_3006_),
    .B(_3004_),
    .Y(\datapath_1.a3 [0])
);

NOR3X1 _13055_ (
    .A(_2611_),
    .B(_2608_),
    .C(_2609_),
    .Y(_2612_)
);

FILL FILL366320x44460 (
);

FILL FILL219640x88920 (
);

FILL FILL_0__14551_ (
);

FILL FILL_0__14131_ (
);

FILL FILL341240x222300 (
);

FILL FILL378480x345800 (
);

FILL FILL_0__9517_ (
);

FILL FILL_0__15756_ (
);

FILL FILL_0__15336_ (
);

AND2X2 _15621_ (
    .A(_4151__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_4573_)
);

AND2X2 _15201_ (
    .A(_4158__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_4159_)
);

FILL FILL_0__10051_ (
);

FILL FILL195320x34580 (
);

AND2X2 _18093_ (
    .A(_6272__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_7008_)
);

FILL FILL_1__17968_ (
);

FILL FILL487920x79040 (
);

AND2X2 _16826_ (
    .A(_5759_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd2 [24])
);

OR2X2 _16406_ (
    .A(_5344_),
    .B(_5345_),
    .Y(_5346_)
);

FILL FILL39520x172900 (
);

FILL FILL_0__9690_ (
);

FILL FILL_0__9270_ (
);

OR2X2 _11961_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [7]),
    .Y(_1799_)
);

DFFSR _11541_ (
    .CLK(clk_bF$buf34),
    .D(_1521_[21]),
    .Q(\datapath_1.regfile_1.regOut[24] [21]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_0__11256_ (
);

OR2X2 _11121_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_1379_)
);

OR2X2 _19298_ (
    .A(_8192_),
    .B(_8193_),
    .Y(_8194_)
);

FILL FILL_0__17902_ (
);

OR2X2 _8748_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_157_)
);

FILL FILL392920x251940 (
);

FILL FILL_1__13048_ (
);

FILL FILL10640x163020 (
);

OR2X2 _12746_ (
    .A(_2267_),
    .B(_2310_),
    .Y(_2311_)
);

OR2X2 _12326_ (
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .Y(_2047_)
);

FILL FILL126920x182780 (
);

FILL FILL_0__13822_ (
);

FILL FILL_0__16294_ (
);

FILL FILL502360x108680 (
);

FILL FILL_1__15614_ (
);

OR2X2 _17784_ (
    .A(_6702_),
    .B(_6703_),
    .Y(_6704_)
);

FILL FILL_0__17079_ (
);

AND2X2 _17364_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_6290_)
);

FILL FILL_0__18860_ (
);

FILL FILL_0__18440_ (
);

OR2X2 _9286_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .B(_464__bF$buf1),
    .Y(_436_)
);

FILL FILL471200x192660 (
);

FILL FILL_1__11114_ (
);

FILL FILL_0__8541_ (
);

FILL FILL_0__10947_ (
);

OR2X2 _10812_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_1213_)
);

FILL FILL_0__10527_ (
);

OR2X2 _18989_ (
    .A(_7888_),
    .B(_7889_),
    .Y(_7890_)
);

AND2X2 _18569_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_7477_)
);

AND2X2 _18149_ (
    .A(_6264__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_7063_)
);

AND2X2 _13284_ (
    .A(_2825_),
    .B(_2826_),
    .Y(_2827_)
);

FILL FILL504640x197600 (
);

FILL FILL485640x153140 (
);

FILL FILL_0__19225_ (
);

AND2X2 _19510_ (
    .A(_8375_),
    .B(_8374_),
    .Y(_8320_[27])
);

FILL FILL_0__14780_ (
);

FILL FILL288040x83980 (
);

DFFSR _14489_ (
    .CLK(clk_bF$buf78),
    .D(_3672_[24]),
    .Q(\datapath_1.Data [24]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _14069_ (
    .A(_3352__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3479_)
);

FILL FILL_1__16572_ (
);

AND2X2 _15850_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_4799_)
);

FILL FILL_0__15565_ (
);

FILL FILL_0__15145_ (
);

AND2X2 _15430_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_4385_)
);

DFFSR _15010_ (
    .CLK(clk_bF$buf12),
    .D(_3936_[29]),
    .Q(\datapath_1.PCJump [29]),
    .R(rst_bF$buf91),
    .S(vdd)
);

FILL FILL_1__17357_ (
);

AND2X2 _16635_ (
    .A(_4200__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_5571_)
);

OR2X2 _16215_ (
    .A(_5157_),
    .B(_5154_),
    .Y(_5158_)
);

FILL FILL_0__11485_ (
);

OR2X2 _11770_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_1718__bF$buf1),
    .Y(_1712_)
);

OR2X2 _11350_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .B(_1520__bF$buf1),
    .Y(_1492_)
);

FILL FILL_0__11065_ (
);

FILL FILL_0__17711_ (
);

OR2X2 _8977_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .B(_332__bF$buf0),
    .Y(_270_)
);

DFFSR _8557_ (
    .CLK(clk_bF$buf51),
    .D(_3_[4]),
    .Q(\datapath_1.regfile_1.regOut[1] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL242440x128440 (
);

FILL FILL_1__10805_ (
);

FILL FILL_1__13697_ (
);

AND2X2 _12975_ (
    .A(_2536_),
    .B(_2534_),
    .Y(_2537_)
);

OR2X2 _12555_ (
    .A(_2138_),
    .B(_2142_),
    .Y(\control_1.next [2])
);

OR2X2 _12135_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_1895_)
);

FILL FILL452200x0 (
);

FILL FILL_0__18916_ (
);

FILL FILL_0__13631_ (
);

FILL FILL_0__13211_ (
);

FILL FILL282720x222300 (
);

FILL FILL_0__14836_ (
);

AND2X2 _14701_ (
    .A(_3853_),
    .B(_3852_),
    .Y(_3804_[24])
);

BUFX2 BUFX2_insert720 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf3 )
);

BUFX2 BUFX2_insert721 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf2 )
);

BUFX2 BUFX2_insert722 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf1 )
);

BUFX2 BUFX2_insert723 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf0 )
);

BUFX2 BUFX2_insert724 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf4 )
);

OR2X2 _17593_ (
    .A(_6515_),
    .B(_6512_),
    .Y(_6516_)
);

BUFX2 BUFX2_insert725 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf3 )
);

BUFX2 BUFX2_insert726 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf2 )
);

AND2X2 _17173_ (
    .A(_4189__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_6101_)
);

FILL FILL32680x44460 (
);

BUFX2 BUFX2_insert727 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf1 )
);

BUFX2 BUFX2_insert728 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf0 )
);

BUFX2 BUFX2_insert729 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf4 )
);

FILL FILL449920x167960 (
);

FILL FILL348840x59280 (
);

DFFSR _9095_ (
    .CLK(clk_bF$buf109),
    .D(_267_[26]),
    .Q(\datapath_1.regfile_1.regOut[5] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

AND2X2 _15906_ (
    .A(_4142__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_4854_)
);

FILL FILL_0__8770_ (
);

DFFSR _10621_ (
    .CLK(clk_bF$buf82),
    .D(_1059_[4]),
    .Q(\datapath_1.regfile_1.regOut[17] [4]),
    .R(rst_bF$buf94),
    .S(vdd)
);

FILL FILL_0__10336_ (
);

OR2X2 _10201_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .B(_926__bF$buf4),
    .Y(_906_)
);

OR2X2 _18798_ (
    .A(_7701_),
    .B(_7700_),
    .Y(_7702_)
);

AND2X2 _18378_ (
    .A(_6211__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_7289_)
);

AND2X2 _13093_ (
    .A(_2306_),
    .B(_2269_),
    .Y(_2648_)
);

FILL FILL_0__19454_ (
);

FILL FILL326040x326040 (
);

FILL FILL_0__9555_ (
);

FILL FILL_0__9135_ (
);

OR2X2 _11826_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_1729_)
);

DFFSR _11406_ (
    .CLK(clk_bF$buf90),
    .D(_1455_[15]),
    .Q(\datapath_1.regfile_1.regOut[23] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL170240x316160 (
);

FILL FILL36480x44460 (
);

OR2X2 _14298_ (
    .A(\datapath_1.ALUResult [19]),
    .B(_3671__bF$buf1),
    .Y(_3645_)
);

FILL FILL_0__15794_ (
);

FILL FILL443840x108680 (
);

FILL FILL174040x237120 (
);

FILL FILL_1__17586_ (
);

FILL FILL_0__16579_ (
);

OR2X2 _16864_ (
    .A(_5793_),
    .B(_5796_),
    .Y(_5797_)
);

FILL FILL_0__16159_ (
);

AND2X2 _16444_ (
    .A(_4177__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_5383_)
);

OR2X2 _16024_ (
    .A(_4962_),
    .B(_4969_),
    .Y(_4970_)
);

FILL FILL_0__11294_ (
);

FILL FILL274360x330980 (
);

FILL FILL_0__17520_ (
);

FILL FILL_0__17100_ (
);

FILL FILL255360x167960 (
);

FILL FILL199880x59280 (
);

AND2X2 _8786_ (
    .A(_182_),
    .B(_181_),
    .Y(_135_[23])
);

FILL FILL25080x172900 (
);

FILL FILL_1__10614_ (
);

FILL FILL16720x14820 (
);

FILL FILL291840x340860 (
);

FILL FILL505400x133380 (
);

OR2X2 _17649_ (
    .A(_6569_),
    .B(_6570_),
    .Y(_6571_)
);

AND2X2 _17229_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_6156_)
);

AND2X2 _12784_ (
    .A(_2343_),
    .B(_2348_),
    .Y(_2349_)
);

FILL FILL_0__12499_ (
);

OR2X2 _12364_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .B(_2048__bF$buf0),
    .Y(_2008_)
);

FILL FILL_0__18725_ (
);

FILL FILL_0__18305_ (
);

FILL FILL_0__13860_ (
);

FILL FILL_0__13440_ (
);

FILL FILL_0__8406_ (
);

AND2X2 _13989_ (
    .A(_3347__bF$buf0),
    .B(\datapath_1.PCJump [12]),
    .Y(_3410_)
);

AND2X2 _13569_ (
    .A(_3067_),
    .B(_3066_),
    .Y(_1_[26])
);

XOR2X1 _13149_ (
    .A(_2696_),
    .B(_2699_),
    .Y(_2700_)
);

FILL FILL_0__14645_ (
);

OR2X2 _14930_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [15]),
    .Y(_3966_)
);

OR2X2 _14510_ (
    .A(IRWrite_bF$buf4),
    .B(\aluControl_1.inst [4]),
    .Y(_3746_)
);

FILL FILL31920x306280 (
);

FILL FILL348840x163020 (
);

FILL FILL370120x281580 (
);

FILL FILL_1__16437_ (
);

FILL FILL367080x232180 (
);

OR2X2 _15715_ (
    .A(_4665_),
    .B(_4664_),
    .Y(_4666_)
);

AND2X2 _10850_ (
    .A(_1238_),
    .B(_1237_),
    .Y(_1191_[23])
);

FILL FILL_0__10565_ (
);

FILL FILL_0__10145_ (
);

AND2X2 _10430_ (
    .A(_1018_),
    .B(_1017_),
    .Y(_993_[12])
);

AND2X2 _10010_ (
    .A(_798_),
    .B(_797_),
    .Y(_795_[1])
);

OR2X2 _18187_ (
    .A(_7100_),
    .B(_7084_),
    .Y(_7101_)
);

FILL FILL384560x242060 (
);

FILL FILL253080x350740 (
);

FILL FILL164920x286520 (
);

FILL FILL280440x59280 (
);

FILL FILL_0__9364_ (
);

OR2X2 _11635_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .B(_1652__bF$buf1),
    .Y(_1642_)
);

OR2X2 _11215_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .B(_1454__bF$buf4),
    .Y(_1422_)
);

FILL FILL270560x360620 (
);

FILL FILL_0__12711_ (
);

FILL FILL384560x108680 (
);

FILL FILL_1__16190_ (
);

FILL FILL455240x69160 (
);

FILL FILL251560x197600 (
);

FILL FILL_0__15183_ (
);

FILL FILL501600x163020 (
);

FILL FILL84360x118560 (
);

FILL FILL_1__14923_ (
);

FILL FILL_0__13916_ (
);

AND2X2 _16673_ (
    .A(_4241__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_5609_)
);

FILL FILL_0__16388_ (
);

OR2X2 _16253_ (
    .A(_5194_),
    .B(_5193_),
    .Y(_5195_)
);

FILL FILL281200x232180 (
);

FILL FILL_1__9525_ (
);

FILL FILL82840x286520 (
);

FILL FILL88160x360620 (
);

OR2X2 _8595_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_75_)
);

FILL FILL_1__10423_ (
);

FILL FILL314640x237120 (
);

AND2X2 _17878_ (
    .A(_6293__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_6796_)
);

AND2X2 _17458_ (
    .A(_6272__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_6383_)
);

AND2X2 _17038_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .Y(_5968_)
);

OR2X2 _12593_ (
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2158_)
);

DFFSR _12173_ (
    .CLK(clk_bF$buf110),
    .D(_1851_[8]),
    .Q(\datapath_1.regfile_1.regOut[29] [8]),
    .R(rst_bF$buf74),
    .S(vdd)
);

FILL FILL_1__19121_ (
);

FILL FILL_0__18954_ (
);

FILL FILL14440x247000 (
);

FILL FILL145160x138320 (
);

FILL FILL350360x316160 (
);

DFFSR _10906_ (
    .CLK(clk_bF$buf83),
    .D(_1191_[31]),
    .Q(\datapath_1.regfile_1.regOut[19] [31]),
    .R(rst_bF$buf81),
    .S(vdd)
);

AND2X2 _13798_ (
    .A(_3089__bF$buf2),
    .B(gnd),
    .Y(_3264_)
);

NAND2X1 _13378_ (
    .A(_2547_),
    .B(_2915_),
    .Y(_2916_)
);

FILL FILL_0__19319_ (
);

FILL FILL_0__14454_ (
);

FILL FILL_0__14034_ (
);

FILL FILL468160x306280 (
);

FILL FILL299440x301340 (
);

FILL FILL82080x301340 (
);

FILL FILL485640x316160 (
);

FILL FILL63080x138320 (
);

OR2X2 _15944_ (
    .A(_4890_),
    .B(_4887_),
    .Y(_4891_)
);

FILL FILL_0__15659_ (
);

AND2X2 _15524_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_4478_)
);

AND2X2 _15104_ (
    .A(_4085_),
    .B(_4029_),
    .Y(\datapath_1.regfile_1.regEn [8])
);

FILL FILL471960x340860 (
);

FILL FILL_0__16600_ (
);

FILL FILL266760x24700 (
);

FILL FILL_0__19492_ (
);

FILL FILL_0__19072_ (
);

OR2X2 _16729_ (
    .A(_5663_),
    .B(_5648_),
    .Y(_5664_)
);

OR2X2 _16309_ (
    .A(_5249_),
    .B(_5250_),
    .Y(_5251_)
);

FILL FILL_0__11999_ (
);

FILL FILL_0__11579_ (
);

AND2X2 _11864_ (
    .A(_1754_),
    .B(_1753_),
    .Y(_1719_[17])
);

AND2X2 _11444_ (
    .A(_1534_),
    .B(_1533_),
    .Y(_1521_[6])
);

DFFSR _11024_ (
    .CLK(clk_bF$buf9),
    .D(_1257_[20]),
    .Q(\datapath_1.regfile_1.regOut[20] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

FILL FILL_0__17805_ (
);

FILL FILL_0__12940_ (
);

FILL FILL51680x232180 (
);

XNOR2X1 _12649_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2214_)
);

OR2X2 _12229_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .B(_1982__bF$buf3),
    .Y(_1938_)
);

FILL FILL41040x192660 (
);

FILL FILL_1__14312_ (
);

FILL FILL_0__13305_ (
);

FILL FILL_0_BUFX2_insert1060 (
);

FILL FILL_0_BUFX2_insert1062 (
);

FILL FILL_0_BUFX2_insert1063 (
);

AND2X2 _16482_ (
    .A(_4172__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_5421_)
);

FILL FILL_0__16197_ (
);

FILL FILL_0_BUFX2_insert1064 (
);

AND2X2 _16062_ (
    .A(_4217__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_5007_)
);

FILL FILL_0_BUFX2_insert1065 (
);

FILL FILL_0_BUFX2_insert1066 (
);

FILL FILL_0_BUFX2_insert1068 (
);

FILL FILL_1__15937_ (
);

FILL FILL278160x321100 (
);

AND2X2 _17687_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_6608_)
);

FILL FILL171760x266760 (
);

FILL FILL319960x34580 (
);

AND2X2 _17267_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_6194_)
);

FILL FILL_1__19350_ (
);

FILL FILL_0__18343_ (
);

OR2X2 _9189_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_391_)
);

FILL FILL_1__11857_ (
);

FILL FILL163400x24700 (
);

AND2X2 _10715_ (
    .A(_1168_),
    .B(_1167_),
    .Y(_1125_[21])
);

FILL FILL252320x133380 (
);

OR2X2 _13187_ (
    .A(_2157__bF$buf3),
    .B(_2735_),
    .Y(_2736_)
);

FILL FILL_1__15690_ (
);

FILL FILL277400x93860 (
);

FILL FILL59280x261820 (
);

FILL FILL461320x93860 (
);

OR2X2 _19413_ (
    .A(_8307_),
    .B(_8304_),
    .Y(_8308_)
);

FILL FILL231800x9880 (
);

FILL FILL_0__14683_ (
);

FILL FILL_0__14263_ (
);

FILL FILL330600x113620 (
);

FILL FILL_0__9649_ (
);

FILL FILL_1__16055_ (
);

FILL FILL_0__15888_ (
);

OR2X2 _15753_ (
    .A(_4695_),
    .B(_4702_),
    .Y(_4703_)
);

FILL FILL_0__15048_ (
);

AND2X2 _15333_ (
    .A(_4210__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_4290_)
);

FILL FILL_0__10183_ (
);

FILL FILL142120x172900 (
);

FILL FILL139080x123500 (
);

FILL FILL9120x143260 (
);

FILL FILL87400x143260 (
);

AND2X2 _16958_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_5889_)
);

AND2X2 _16538_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_5476_)
);

OR2X2 _16118_ (
    .A(_5059_),
    .B(_5062_),
    .Y(_5063_)
);

FILL FILL_0__11388_ (
);

DFFSR _11673_ (
    .CLK(clk_bF$buf96),
    .D(_1587_[24]),
    .Q(\datapath_1.regfile_1.regOut[25] [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL_1__18201_ (
);

OR2X2 _11253_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_1447_)
);

FILL FILL38760x330980 (
);

FILL FILL_1__10708_ (
);

AND2X2 _9821_ (
    .A(_712_),
    .B(_711_),
    .Y(_663_[24])
);

AND2X2 _9401_ (
    .A(_492_),
    .B(_491_),
    .Y(_465_[13])
);

OR2X2 _12878_ (
    .A(_2441_),
    .B(_2442_),
    .Y(_2443_)
);

NAND3X1 _12458_ (
    .A(_2051_),
    .B(_2049_),
    .C(\aluControl_1.inst [2]),
    .Y(_2052_)
);

DFFSR _12038_ (
    .CLK(clk_bF$buf18),
    .D(_1785_[2]),
    .Q(\datapath_1.regfile_1.regOut[28] [2]),
    .R(rst_bF$buf107),
    .S(vdd)
);

FILL FILL_1__14961_ (
);

FILL FILL_0__18819_ (
);

FILL FILL287280x118560 (
);

FILL FILL_0__13954_ (
);

FILL FILL374680x123500 (
);

FILL FILL_0__13534_ (
);

FILL FILL_0__13114_ (
);

FILL FILL231040x153140 (
);

FILL FILL502360x29640 (
);

OR2X2 _16291_ (
    .A(_5231_),
    .B(_5232_),
    .Y(_5233_)
);

DFFSR _14604_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[10]),
    .Q(\datapath_1.PCJump [12]),
    .R(rst_bF$buf100),
    .S(vdd)
);

OR2X2 _17496_ (
    .A(_6416_),
    .B(_6419_),
    .Y(_6420_)
);

AND2X2 _17076_ (
    .A(_4210__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_6006_)
);

FILL FILL_0__18992_ (
);

FILL FILL_0__18572_ (
);

FILL FILL_0__18152_ (
);

OR2X2 _15809_ (
    .A(_4757_),
    .B(_4754_),
    .Y(_4758_)
);

FILL FILL268280x0 (
);

FILL FILL_0__8673_ (
);

FILL FILL_0__10659_ (
);

OR2X2 _10944_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_1281_)
);

OR2X2 _10524_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_1061_)
);

DFFSR _10104_ (
    .CLK(clk_bF$buf71),
    .D(_795_[3]),
    .Q(\datapath_1.regfile_1.regOut[13] [3]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL_0__11600_ (
);

FILL FILL_0__19357_ (
);

AND2X2 _19222_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_8120_)
);

FILL FILL251560x34580 (
);

FILL FILL_0__14072_ (
);

FILL FILL25840x54340 (
);

FILL FILL_0__9038_ (
);

AND2X2 _11729_ (
    .A(_1684_),
    .B(_1683_),
    .Y(_1653_[15])
);

AND2X2 _11309_ (
    .A(_1464_),
    .B(_1463_),
    .Y(_1455_[4])
);

FILL FILL161880x69160 (
);

FILL FILL110200x316160 (
);

FILL FILL179360x227240 (
);

FILL FILL_0__12805_ (
);

FILL FILL38000x296400 (
);

OR2X2 _15982_ (
    .A(_4927_),
    .B(_4928_),
    .Y(_4929_)
);

FILL FILL_0__15697_ (
);

FILL FILL_0__15277_ (
);

AND2X2 _15562_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_4515_)
);

NAND2X1 _15142_ (
    .A(\datapath_1.a3 [4]),
    .B(_4079_),
    .Y(_4110_)
);

FILL FILL458280x321100 (
);

FILL FILL22040x69160 (
);

FILL FILL278920x34580 (
);

FILL FILL462840x34580 (
);

FILL FILL283480x148200 (
);

AND2X2 _16767_ (
    .A(_4189__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_5701_)
);

AND2X2 _16347_ (
    .A(_4177__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_5288_)
);

FILL FILL255360x34580 (
);

FILL FILL_1__18850_ (
);

OR2X2 _11482_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .B(_1586__bF$buf0),
    .Y(_1560_)
);

FILL FILL_0__11197_ (
);

OR2X2 _11062_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_1388__bF$buf4),
    .Y(_1340_)
);

FILL FILL_1__9619_ (
);

FILL FILL_0__17843_ (
);

FILL FILL_0__17423_ (
);

FILL FILL15200x321100 (
);

DFFSR _8689_ (
    .CLK(clk_bF$buf48),
    .D(_69_[7]),
    .Q(\datapath_1.regfile_1.regOut[2] [7]),
    .R(rst_bF$buf21),
    .S(vdd)
);

FILL FILL165680x69160 (
);

OR2X2 _9630_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_605_)
);

DFFSR _9210_ (
    .CLK(clk_bF$buf106),
    .D(_333_[12]),
    .Q(\datapath_1.regfile_1.regOut[6] [12]),
    .R(rst_bF$buf0),
    .S(vdd)
);

INVX1 _12687_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .Y(_2252_)
);

FILL FILL_1__19215_ (
);

OR2X2 _12267_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_1963_)
);

FILL FILL505400x247000 (
);

FILL FILL_1__14770_ (
);

AND2X2 _18913_ (
    .A(_6221__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_7815_)
);

FILL FILL_0__18208_ (
);

FILL FILL_0__13763_ (
);

FILL FILL_0__8729_ (
);

FILL FILL_1__15555_ (
);

FILL FILL_0__14968_ (
);

FILL FILL313880x370500 (
);

AND2X2 _14833_ (
    .A(_3921_),
    .B(_3920_),
    .Y(_3870_[25])
);

FILL FILL_0__14128_ (
);

AND2X2 _14413_ (
    .A(_3701_),
    .B(_3700_),
    .Y(_3672_[14])
);

FILL FILL145920x39520 (
);

FILL FILL_1__11475_ (
);

AND2X2 _15618_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_4570_)
);

FILL FILL_0__10468_ (
);

DFFSR _10753_ (
    .CLK(clk_bF$buf18),
    .D(_1125_[7]),
    .Q(\datapath_1.regfile_1.regOut[18] [7]),
    .R(rst_bF$buf107),
    .S(vdd)
);

OR2X2 _10333_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .B(_992__bF$buf0),
    .Y(_974_)
);

OR2X2 _19451_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_8336_)
);

FILL FILL_0__19166_ (
);

OR2X2 _19031_ (
    .A(_7924_),
    .B(_7931_),
    .Y(_7932_)
);

FILL FILL441560x14820 (
);

OR2X2 _8901_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_239_)
);

FILL FILL298680x113620 (
);

FILL FILL_0__9267_ (
);

OR2X2 _11958_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_1797_)
);

DFFSR _11538_ (
    .CLK(clk_bF$buf61),
    .D(_1521_[18]),
    .Q(\datapath_1.regfile_1.regOut[24] [18]),
    .R(rst_bF$buf11),
    .S(vdd)
);

OR2X2 _11118_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_1377_)
);

FILL FILL217360x64220 (
);

FILL FILL_0__12614_ (
);

FILL FILL207480x311220 (
);

FILL FILL348080x83980 (
);

OR2X2 _15791_ (
    .A(_4740_),
    .B(_4737_),
    .Y(_4741_)
);

AND2X2 _15371_ (
    .A(_4239__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_4327_)
);

FILL FILL140600x365560 (
);

FILL FILL44840x24700 (
);

FILL FILL104880x177840 (
);

AND2X2 _16996_ (
    .A(_4160__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_5927_)
);

OR2X2 _16576_ (
    .A(_5512_),
    .B(_5511_),
    .Y(_5513_)
);

FILL FILL144400x286520 (
);

OR2X2 _16156_ (
    .A(_5099_),
    .B(_5098_),
    .Y(_5100_)
);

DFFSR _11291_ (
    .CLK(clk_bF$buf64),
    .D(_1389_[29]),
    .Q(\datapath_1.regfile_1.regOut[22] [29]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL_1__9428_ (
);

AND2X2 _8498_ (
    .A(_30_),
    .B(_29_),
    .Y(_3_[13])
);

FILL FILL476520x158080 (
);

FILL FILL465120x29640 (
);

NAND2X1 _12496_ (
    .A(_2097_),
    .B(_2096_),
    .Y(_2098_)
);

OR2X2 _12076_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .B(_1916__bF$buf2),
    .Y(_1856_)
);

FILL FILL_0__18857_ (
);

AND2X2 _18722_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_7627_)
);

FILL FILL_0__18437_ (
);

AND2X2 _18302_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_7214_)
);

FILL FILL_0__18017_ (
);

FILL FILL_0__13152_ (
);

FILL FILL_0__8538_ (
);

OR2X2 _10809_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_1211_)
);

FILL FILL102600x148200 (
);

FILL FILL62320x286520 (
);

FILL FILL385320x360620 (
);

FILL FILL215080x88920 (
);

FILL FILL499320x108680 (
);

AND2X2 _19507_ (
    .A(_8373_),
    .B(_8372_),
    .Y(_8320_[26])
);

FILL FILL114000x64220 (
);

OR2X2 _14642_ (
    .A(vdd),
    .B(\datapath_1.a [5]),
    .Y(_3814_)
);

OR2X2 _14222_ (
    .A(\datapath_1.Data [26]),
    .B(_3605__bF$buf0),
    .Y(_3593_)
);

FILL FILL_0__18190_ (
);

FILL FILL449920x88920 (
);

FILL FILL425600x316160 (
);

OR2X2 _15847_ (
    .A(_4795_),
    .B(_4792_),
    .Y(_4796_)
);

AND2X2 _15427_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_4382_)
);

DFFSR _15007_ (
    .CLK(clk_bF$buf77),
    .D(_3936_[26]),
    .Q(\datapath_1.mux_iord.din0 [26]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL_0__10697_ (
);

AND2X2 _10982_ (
    .A(_1306_),
    .B(_1305_),
    .Y(_1257_[24])
);

AND2X2 _10562_ (
    .A(_1086_),
    .B(_1085_),
    .Y(_1059_[13])
);

FILL FILL_0__10277_ (
);

FILL FILL389120x44460 (
);

AND2X2 _10142_ (
    .A(_866_),
    .B(_865_),
    .Y(_861_[2])
);

FILL FILL_0__16923_ (
);

FILL FILL_0__16503_ (
);

FILL FILL408880x59280 (
);

FILL FILL20520x148200 (
);

FILL FILL_0__19395_ (
);

OR2X2 _19260_ (
    .A(_8156_),
    .B(_8142_),
    .Y(_8157_)
);

FILL FILL483360x79040 (
);

DFFSR _8710_ (
    .CLK(clk_bF$buf72),
    .D(_69_[28]),
    .Q(\datapath_1.regfile_1.regOut[2] [28]),
    .R(rst_bF$buf89),
    .S(vdd)
);

OR2X2 _11767_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .B(_1718__bF$buf2),
    .Y(_1710_)
);

FILL FILL_1__18715_ (
);

OR2X2 _11347_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .B(_1520__bF$buf0),
    .Y(_1490_)
);

FILL FILL159600x251940 (
);

FILL FILL_1__13430_ (
);

FILL FILL435480x0 (
);

FILL FILL_0__12003_ (
);

FILL FILL296400x0 (
);

INVX1 _15180_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_4138_)
);

OR2X2 _9915_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_755_)
);

AND2X2 _13913_ (
    .A(_3343_),
    .B(ALUSrcB[0]),
    .Y(_3344_)
);

FILL FILL_0__13628_ (
);

FILL FILL392160x113620 (
);

OR2X2 _16385_ (
    .A(_5321_),
    .B(_5324_),
    .Y(_5325_)
);

FILL FILL200640x103740 (
);

FILL FILL_1__9237_ (
);

FILL FILL_0__17461_ (
);

FILL FILL_0__17041_ (
);

FILL FILL110960x34580 (
);

FILL FILL_1__10555_ (
);

BUFX2 BUFX2_insert690 (
    .A(_6238_),
    .Y(_6238__bF$buf4)
);

BUFX2 BUFX2_insert691 (
    .A(_6238_),
    .Y(_6238__bF$buf3)
);

BUFX2 BUFX2_insert692 (
    .A(_6238_),
    .Y(_6238__bF$buf2)
);

BUFX2 BUFX2_insert693 (
    .A(_6238_),
    .Y(_6238__bF$buf1)
);

BUFX2 BUFX2_insert694 (
    .A(_6238_),
    .Y(_6238__bF$buf0)
);

BUFX2 BUFX2_insert695 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf4 )
);

BUFX2 BUFX2_insert696 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf3 )
);

BUFX2 BUFX2_insert697 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf2 )
);

BUFX2 BUFX2_insert698 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf1 )
);

BUFX2 BUFX2_insert699 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf0 )
);

FILL FILL_0__18666_ (
);

AND2X2 _18951_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_7853_)
);

FILL FILL_0__18246_ (
);

OR2X2 _18531_ (
    .A(_7430_),
    .B(_7438_),
    .Y(_7439_)
);

AND2X2 _18111_ (
    .A(_6262__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_7026_)
);

FILL FILL_0__13381_ (
);

FILL FILL504640x108680 (
);

FILL FILL90440x93860 (
);

FILL FILL307800x370500 (
);

DFFSR _10618_ (
    .CLK(clk_bF$buf85),
    .D(_1059_[1]),
    .Q(\datapath_1.regfile_1.regOut[17] [1]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL_1__15173_ (
);

OR2X2 _19316_ (
    .A(_8208_),
    .B(_8211_),
    .Y(_8212_)
);

DFFSR _14871_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[19]),
    .Q(_2_[19]),
    .R(rst_bF$buf61),
    .S(vdd)
);

FILL FILL_0__14586_ (
);

OR2X2 _14451_ (
    .A(memoryOutData[27]),
    .B(_3737__bF$buf0),
    .Y(_3727_)
);

AND2X2 _14031_ (
    .A(_3347__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3446_)
);

FILL FILL_1__16378_ (
);

OR2X2 _15656_ (
    .A(_4607_),
    .B(_4600_),
    .Y(_4608_)
);

OR2X2 _15236_ (
    .A(_4164_),
    .B(_4193_),
    .Y(_4194_)
);

OR2X2 _10791_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_1199_)
);

DFFSR _10371_ (
    .CLK(clk_bF$buf75),
    .D(_927_[12]),
    .Q(\datapath_1.regfile_1.regOut[15] [12]),
    .R(rst_bF$buf27),
    .S(vdd)
);

FILL FILL_0__10086_ (
);

FILL FILL487920x153140 (
);

FILL FILL_1__8508_ (
);

FILL FILL_0__16312_ (
);

FILL FILL56240x271700 (
);

AND2X2 _11996_ (
    .A(_1822_),
    .B(_1821_),
    .Y(_1785_[18])
);

FILL FILL301720x311220 (
);

AND2X2 _11576_ (
    .A(_1602_),
    .B(_1601_),
    .Y(_1587_[7])
);

DFFSR _11156_ (
    .CLK(clk_bF$buf87),
    .D(_1323_[23]),
    .Q(\datapath_1.regfile_1.regOut[21] [23]),
    .R(rst_bF$buf54),
    .S(vdd)
);

FILL FILL392160x340860 (
);

FILL FILL_0__17937_ (
);

FILL FILL_0__17517_ (
);

AND2X2 _17802_ (
    .A(_6326__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_6721_)
);

FILL FILL_0__12652_ (
);

FILL FILL174040x88920 (
);

DFFSR _9724_ (
    .CLK(clk_bF$buf33),
    .D(_597_[10]),
    .Q(\datapath_1.regfile_1.regOut[10] [10]),
    .R(rst_bF$buf56),
    .S(vdd)
);

OR2X2 _9304_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .B(_464__bF$buf0),
    .Y(_448_)
);

FILL FILL104880x247000 (
);

OR2X2 _13722_ (
    .A(_3198_),
    .B(_3197_),
    .Y(_3199_)
);

FILL FILL_0__13017_ (
);

XOR2X1 _13302_ (
    .A(_2425_),
    .B(_2415_),
    .Y(_2844_)
);

AND2X2 _16194_ (
    .A(_4130__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_5137_)
);

FILL FILL500840x138320 (
);

FILL FILL244720x128440 (
);

FILL FILL_0__17690_ (
);

FILL FILL_0__17270_ (
);

OR2X2 _14927_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [14]),
    .Y(_3964_)
);

OR2X2 _14507_ (
    .A(IRWrite_bF$buf4),
    .B(\aluControl_1.inst [3]),
    .Y(_3744_)
);

FILL FILL449160x163020 (
);

OR2X2 _17399_ (
    .A(_6322_),
    .B(_6324_),
    .Y(_6325_)
);

FILL FILL320720x29640 (
);

FILL FILL344280x59280 (
);

FILL FILL_0__18895_ (
);

AND2X2 _18760_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_7665_)
);

FILL FILL_0__18475_ (
);

OR2X2 _18340_ (
    .A(_7249_),
    .B(_7250_),
    .Y(_7251_)
);

FILL FILL_0__13190_ (
);

FILL FILL_1__11569_ (
);

FILL FILL_0__8996_ (
);

AND2X2 _10847_ (
    .A(_1236_),
    .B(_1235_),
    .Y(_1191_[22])
);

AND2X2 _10427_ (
    .A(_1016_),
    .B(_1015_),
    .Y(_993_[11])
);

AND2X2 _10007_ (
    .A(_796_),
    .B(_859_),
    .Y(_795_[0])
);

DFFSR _19545_ (
    .CLK(clk_bF$buf91),
    .D(_8320_[22]),
    .Q(\datapath_1.regfile_1.regOut[0] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

AND2X2 _19125_ (
    .A(_6264__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_8024_)
);

AND2X2 _14680_ (
    .A(_3839_),
    .B(_3838_),
    .Y(_3804_[17])
);

FILL FILL_0__14395_ (
);

AND2X2 _14260_ (
    .A(_3619_),
    .B(_3618_),
    .Y(_3606_[6])
);

FILL FILL489440x123500 (
);

FILL FILL79040x365560 (
);

FILL FILL11400x79040 (
);

AND2X2 _15885_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_4833_)
);

AND2X2 _15465_ (
    .A(_4241__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_4420_)
);

AND2X2 _15045_ (
    .A(_4032_),
    .B(_4033_),
    .Y(_4034_)
);

FILL FILL91960x34580 (
);

OR2X2 _10180_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .B(_926__bF$buf1),
    .Y(_892_)
);

FILL FILL_0__16961_ (
);

FILL FILL_0__16541_ (
);

FILL FILL155040x306280 (
);

FILL FILL_1__18333_ (
);

OR2X2 _11385_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_1515_)
);

OR2X2 _17611_ (
    .A(_6531_),
    .B(_6532_),
    .Y(_6533_)
);

FILL FILL_0__17326_ (
);

FILL FILL_0__12881_ (
);

FILL FILL_0__12461_ (
);

FILL FILL340480x291460 (
);

FILL FILL409640x256880 (
);

FILL FILL145160x251940 (
);

AND2X2 _9953_ (
    .A(_780_),
    .B(_779_),
    .Y(_729_[25])
);

AND2X2 _9533_ (
    .A(_560_),
    .B(_559_),
    .Y(_531_[14])
);

AND2X2 _9113_ (
    .A(_340_),
    .B(_339_),
    .Y(_333_[3])
);

FILL FILL_1__14673_ (
);

OR2X2 _18816_ (
    .A(_7718_),
    .B(_7719_),
    .Y(_7720_)
);

FILL FILL_0_BUFX2_insert330 (
);

FILL FILL_0_BUFX2_insert331 (
);

FILL FILL_0_BUFX2_insert333 (
);

OR2X2 _13951_ (
    .A(_3377_),
    .B(_3376_),
    .Y(_3378_)
);

FILL FILL_0__13666_ (
);

FILL FILL_0__13246_ (
);

FILL FILL_0_BUFX2_insert335 (
);

OR2X2 _13531_ (
    .A(IorD_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [14]),
    .Y(_3042_)
);

INVX1 _13111_ (
    .A(_2664_),
    .Y(\datapath_1.ALUResult [20])
);

FILL FILL12920x88920 (
);

FILL FILL_0_BUFX2_insert337 (
);

FILL FILL276640x330980 (
);

FILL FILL_0_BUFX2_insert339 (
);

FILL FILL39520x14820 (
);

FILL FILL_1__15038_ (
);

FILL FILL452200x59280 (
);

DFFSR _14736_ (
    .CLK(clk_bF$buf4),
    .D(_3804_[13]),
    .Q(\datapath_1.a [13]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _14316_ (
    .A(\datapath_1.ALUResult [25]),
    .B(_3671__bF$buf3),
    .Y(_3657_)
);

FILL FILL202920x217360 (
);

FILL FILL63080x251940 (
);

FILL FILL_0__15812_ (
);

FILL FILL_1__19291_ (
);

FILL FILL_0__18284_ (
);

OR2X2 _10656_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_1129_)
);

FILL FILL16720x88920 (
);

DFFSR _10236_ (
    .CLK(clk_bF$buf49),
    .D(_861_[6]),
    .Q(\datapath_1.regfile_1.regOut[14] [6]),
    .R(rst_bF$buf106),
    .S(vdd)
);

FILL FILL454480x54340 (
);

FILL FILL_0__11732_ (
);

FILL FILL_0__19489_ (
);

OR2X2 _19354_ (
    .A(_8248_),
    .B(_8249_),
    .Y(_8250_)
);

AND2X2 _8804_ (
    .A(_194_),
    .B(_193_),
    .Y(_135_[29])
);

FILL FILL251560x108680 (
);

FILL FILL_1__13944_ (
);

FILL FILL_1__13524_ (
);

FILL FILL46360x158080 (
);

FILL FILL369360x232180 (
);

NAND2X1 _12802_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(_2352_),
    .Y(_2367_)
);

FILL FILL_0__12517_ (
);

AND2X2 _15694_ (
    .A(_4130__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_4645_)
);

OR2X2 _15274_ (
    .A(_4229_),
    .B(_4231_),
    .Y(_4232_)
);

FILL FILL304000x242060 (
);

AND2X2 _16899_ (
    .A(_4154__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_5831_)
);

OR2X2 _16479_ (
    .A(_5417_),
    .B(_5416_),
    .Y(_5418_)
);

FILL FILL272840x360620 (
);

AND2X2 _16059_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_5004_)
);

FILL FILL_1__18982_ (
);

FILL FILL166440x83980 (
);

OR2X2 _11194_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .B(_1454__bF$buf3),
    .Y(_1408_)
);

FILL FILL386840x108680 (
);

FILL FILL_0__17975_ (
);

FILL FILL253840x197600 (
);

FILL FILL_0__17555_ (
);

AND2X2 _17840_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_6759_)
);

OR2X2 _17420_ (
    .A(_6344_),
    .B(_6343_),
    .Y(_6345_)
);

FILL FILL_0__17135_ (
);

FILL FILL259160x271700 (
);

OR2X2 _17000_ (
    .A(_5923_),
    .B(_5930_),
    .Y(_5931_)
);

FILL FILL_0__12270_ (
);

OR2X2 _9762_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_673_)
);

DFFSR _9342_ (
    .CLK(clk_bF$buf48),
    .D(_399_[15]),
    .Q(\datapath_1.regfile_1.regOut[7] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

OR2X2 _12399_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_2031_)
);

FILL FILL263720x14820 (
);

OR2X2 _18625_ (
    .A(_7528_),
    .B(_7531_),
    .Y(_7532_)
);

OR2X2 _18205_ (
    .A(_7110_),
    .B(_7117_),
    .Y(_7118_)
);

FILL FILL496280x103740 (
);

FILL FILL_0__13895_ (
);

FILL FILL_0__13475_ (
);

AND2X2 _13760_ (
    .A(_3084__bF$buf4),
    .B(\datapath_1.PCJump [24]),
    .Y(_3231_)
);

FILL FILL_0__13055_ (
);

NAND2X1 _13340_ (
    .A(_2524_),
    .B(_2879_),
    .Y(_2880_)
);

FILL FILL143640x217360 (
);

FILL FILL_0__9802_ (
);

AND2X2 _14965_ (
    .A(_3989_),
    .B(_3988_),
    .Y(_3936_[26])
);

AND2X2 _14545_ (
    .A(_3769_),
    .B(_3768_),
    .Y(_3738_[15])
);

AND2X2 _14125_ (
    .A(_3352__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3527_)
);

FILL FILL53200x103740 (
);

FILL FILL321480x330980 (
);

FILL FILL_0__15621_ (
);

FILL FILL180120x44460 (
);

FILL FILL234080x370500 (
);

FILL FILL264480x281580 (
);

FILL FILL_1__17833_ (
);

DFFSR _10885_ (
    .CLK(clk_bF$buf49),
    .D(_1191_[10]),
    .Q(\datapath_1.regfile_1.regOut[19] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

OR2X2 _10465_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .B(_1058__bF$buf2),
    .Y(_1042_)
);

OR2X2 _10045_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .B(_860__bF$buf0),
    .Y(_822_)
);

FILL FILL270560x222300 (
);

FILL FILL348080x118560 (
);

FILL FILL_0__16406_ (
);

FILL FILL_0__11961_ (
);

FILL FILL207480x19760 (
);

FILL FILL_0__19298_ (
);

OR2X2 _19163_ (
    .A(_8029_),
    .B(_8061_),
    .Y(_8062_)
);

OR2X2 _8613_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_87_)
);

FILL FILL_0__9399_ (
);

FILL FILL65360x138320 (
);

FILL FILL_0__12746_ (
);

OR2X2 _12611_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(_2175_),
    .Y(_2176_)
);

FILL FILL_0__12326_ (
);

AND2X2 _15083_ (
    .A(_4068_),
    .B(_4029_),
    .Y(\datapath_1.regfile_1.regEn [4])
);

AND2X2 _9818_ (
    .A(_710_),
    .B(_709_),
    .Y(_663_[23])
);

FILL FILL473480x24700 (
);

FILL FILL418760x19760 (
);

FILL FILL92720x49400 (
);

INVX2 _13816_ (
    .A(ALUSrcA_bF$buf1),
    .Y(_3342_)
);

FILL FILL493240x39520 (
);

OR2X2 _16288_ (
    .A(_5226_),
    .B(_5229_),
    .Y(_5230_)
);

FILL FILL386080x286520 (
);

FILL FILL_0__17784_ (
);

FILL FILL_0__17364_ (
);

FILL FILL53960x232180 (
);

FILL FILL450680x98800 (
);

DFFSR _9991_ (
    .CLK(clk_bF$buf99),
    .D(_729_[19]),
    .Q(\datapath_1.regfile_1.regOut[12] [19]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9571_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .B(_596__bF$buf3),
    .Y(_586_)
);

OR2X2 _9151_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .B(_398__bF$buf3),
    .Y(_366_)
);

FILL FILL43320x192660 (
);

FILL FILL285000x202540 (
);

FILL FILL_1__19156_ (
);

FILL FILL_0__18989_ (
);

FILL FILL_0_BUFX2_insert710 (
);

OR2X2 _18854_ (
    .A(_7756_),
    .B(_7753_),
    .Y(_7757_)
);

FILL FILL_0_BUFX2_insert711 (
);

OR2X2 _18434_ (
    .A(_7343_),
    .B(_7342_),
    .Y(_7344_)
);

OR2X2 _18014_ (
    .A(_6928_),
    .B(_6929_),
    .Y(_6930_)
);

FILL FILL_0_BUFX2_insert713 (
);

FILL FILL_0_BUFX2_insert715 (
);

FILL FILL_0_BUFX2_insert717 (
);

FILL FILL_0_BUFX2_insert719 (
);

FILL FILL383040x182780 (
);

FILL FILL_1__15496_ (
);

AND2X2 _19219_ (
    .A(_6250__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_8117_)
);

OR2X2 _14774_ (
    .A(vdd),
    .B(_2_[6]),
    .Y(_3882_)
);

FILL FILL_0__14069_ (
);

DFFSR _14354_ (
    .CLK(clk_bF$buf77),
    .D(_3606_[18]),
    .Q(ALUOut[18]),
    .R(rst_bF$buf63),
    .S(vdd)
);

FILL FILL29640x286520 (
);

FILL FILL_0__15430_ (
);

FILL FILL_1__13809_ (
);

FILL FILL196840x350740 (
);

FILL FILL297160x237120 (
);

FILL FILL254600x133380 (
);

OR2X2 _15979_ (
    .A(_4924_),
    .B(_4925_),
    .Y(_4926_)
);

OR2X2 _15559_ (
    .A(_4511_),
    .B(_4510_),
    .Y(_4512_)
);

AOI21X1 _15139_ (
    .A(_4002_),
    .B(_4020_),
    .C(_4107_),
    .Y(_4108_)
);

AND2X2 _10694_ (
    .A(_1154_),
    .B(_1153_),
    .Y(_1125_[14])
);

AND2X2 _10274_ (
    .A(_934_),
    .B(_933_),
    .Y(_927_[3])
);

FILL FILL_0__16635_ (
);

OR2X2 _16920_ (
    .A(_5844_),
    .B(_5851_),
    .Y(_5852_)
);

AND2X2 _16500_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_5439_)
);

FILL FILL209000x256880 (
);

FILL FILL_0__11770_ (
);

AND2X2 _19392_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_8287_)
);

DFFSR _8842_ (
    .CLK(clk_bF$buf10),
    .D(_135_[31]),
    .Q(\datapath_1.regfile_1.regOut[3] [31]),
    .R(rst_bF$buf44),
    .S(vdd)
);

BUFX2 _8422_ (
    .A(_1_[30]),
    .Y(memoryAddress[30])
);

OR2X2 _11899_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .B(_1784__bF$buf2),
    .Y(_1778_)
);

OR2X2 _11479_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .B(_1586__bF$buf3),
    .Y(_1558_)
);

OR2X2 _11059_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .B(_1388__bF$buf3),
    .Y(_1338_)
);

FILL FILL_1__18007_ (
);

FILL FILL_1__13562_ (
);

FILL FILL332120x340860 (
);

AND2X2 _17705_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_6626_)
);

FILL FILL212040x34580 (
);

OR2X2 _12840_ (
    .A(_2404_),
    .B(_2400_),
    .Y(_2405_)
);

FILL FILL_0__12135_ (
);

OR2X2 _12420_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_2045_)
);

FILL FILL505400x360620 (
);

OR2X2 _12000_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_1825_)
);

FILL FILL249280x158080 (
);

OR2X2 _9627_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_603_)
);

DFFSR _9207_ (
    .CLK(clk_bF$buf24),
    .D(_333_[9]),
    .Q(\datapath_1.regfile_1.regOut[6] [9]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL319200x19760 (
);

FILL FILL504640x79040 (
);

FILL FILL275120x291460 (
);

OR2X2 _13625_ (
    .A(_3115_),
    .B(_3112_),
    .Y(\datapath_1.mux_pcsrc.dout [4])
);

XOR2X1 _13205_ (
    .A(_2418_),
    .B(_2732_),
    .Y(_2753_)
);

AND2X2 _16097_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_5042_)
);

FILL FILL_0__14701_ (
);

FILL FILL_1__9369_ (
);

FILL FILL_0__17593_ (
);

FILL FILL359480x113620 (
);

FILL FILL_1__10687_ (
);

AND2X2 _9380_ (
    .A(_478_),
    .B(_477_),
    .Y(_465_[6])
);

FILL FILL_0__15906_ (
);

FILL FILL289560x118560 (
);

FILL FILL376960x123500 (
);

INVX1 _18663_ (
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_7569_)
);

FILL FILL_0__18378_ (
);

OR2X2 _18243_ (
    .A(_7155_),
    .B(_7152_),
    .Y(_7156_)
);

FILL FILL_0__13093_ (
);

FILL FILL_0__8479_ (
);

FILL FILL_0__9840_ (
);

FILL FILL_0__9420_ (
);

FILL FILL_0__11826_ (
);

OR2X2 _19448_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [7]),
    .Y(_8334_)
);

AND2X2 _19028_ (
    .A(_6328__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_7929_)
);

OR2X2 _14583_ (
    .A(memoryOutData[28]),
    .B(_3803__bF$buf1),
    .Y(_3795_)
);

AND2X2 _14163_ (
    .A(_3553_),
    .B(_3552_),
    .Y(\datapath_1.mux_wd3.dout [6])
);

FILL FILL21280x54340 (
);

FILL FILL93480x370500 (
);

FILL FILL228000x370500 (
);

FILL FILL384560x335920 (
);

FILL FILL_1_BUFX2_insert260 (
);

FILL FILL_1_BUFX2_insert262 (
);

FILL FILL_1_BUFX2_insert264 (
);

FILL FILL325280x321100 (
);

FILL FILL442320x118560 (
);

FILL FILL481840x34580 (
);

AND2X2 _15788_ (
    .A(_4167__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_4738_)
);

OR2X2 _15368_ (
    .A(_4320_),
    .B(_4323_),
    .Y(_4324_)
);

FILL FILL_1__17451_ (
);

OR2X2 _10083_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_847_)
);

FILL FILL_0__16444_ (
);

FILL FILL_0__16024_ (
);

AND2X2 _8651_ (
    .A(_112_),
    .B(_111_),
    .Y(_69_[21])
);

FILL FILL184680x69160 (
);

FILL FILL437760x237120 (
);

FILL FILL_1__18656_ (
);

DFFSR _11288_ (
    .CLK(clk_bF$buf89),
    .D(_1389_[26]),
    .Q(\datapath_1.regfile_1.regOut[22] [26]),
    .R(rst_bF$buf24),
    .S(vdd)
);

FILL FILL25080x54340 (
);

FILL FILL281960x227240 (
);

FILL FILL_0__17649_ (
);

AND2X2 _17934_ (
    .A(_6216__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_6851_)
);

FILL FILL_0__17229_ (
);

AND2X2 _17514_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_6438_)
);

FILL FILL_0__12784_ (
);

DFFSR _9856_ (
    .CLK(clk_bF$buf13),
    .D(_663_[13]),
    .Q(\datapath_1.regfile_1.regOut[11] [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

OR2X2 _9436_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .B(_530__bF$buf4),
    .Y(_516_)
);

OR2X2 _9016_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_332__bF$buf1),
    .Y(_296_)
);

AND2X2 _18719_ (
    .A(_6255__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_7624_)
);

FILL FILL_0__13989_ (
);

AND2X2 _13854_ (
    .A(_3302_),
    .B(_3301_),
    .Y(\datapath_1.alu_1.ALUInA [12])
);

FILL FILL_0__13569_ (
);

FILL FILL278160x34580 (
);

NAND3X1 _13434_ (
    .A(_2383_),
    .B(_2500_),
    .C(_2967_),
    .Y(_2968_)
);

AND2X2 _13014_ (
    .A(_2572_),
    .B(_2331_),
    .Y(_2573_)
);

FILL FILL_0__14930_ (
);

FILL FILL_0__14510_ (
);

FILL FILL164920x39520 (
);

FILL FILL188480x69160 (
);

OR2X2 _14639_ (
    .A(vdd),
    .B(\datapath_1.a [4]),
    .Y(_3812_)
);

OR2X2 _14219_ (
    .A(\datapath_1.Data [25]),
    .B(_3605__bF$buf1),
    .Y(_3591_)
);

FILL FILL339720x49400 (
);

FILL FILL_1__16302_ (
);

FILL FILL440040x301340 (
);

FILL FILL_0__10850_ (
);

FILL FILL_0__10430_ (
);

OR2X2 _18892_ (
    .A(_7794_),
    .B(_7793_),
    .Y(_7795_)
);

AND2X2 _18472_ (
    .A(_6206__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_7381_)
);

AND2X2 _18052_ (
    .A(_6302__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_6968_)
);

FILL FILL406600x88920 (
);

AND2X2 _10979_ (
    .A(_1304_),
    .B(_1303_),
    .Y(_1257_[23])
);

AND2X2 _10559_ (
    .A(_1084_),
    .B(_1083_),
    .Y(_1059_[12])
);

AND2X2 _10139_ (
    .A(_864_),
    .B(_863_),
    .Y(_861_[1])
);

FILL FILL_1__12642_ (
);

DFFSR _11920_ (
    .CLK(clk_bF$buf103),
    .D(_1719_[13]),
    .Q(\datapath_1.regfile_1.regOut[27] [13]),
    .R(rst_bF$buf32),
    .S(vdd)
);

OR2X2 _11500_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .B(_1586__bF$buf0),
    .Y(_1572_)
);

FILL FILL_0__11215_ (
);

OR2X2 _19257_ (
    .A(_8152_),
    .B(_8153_),
    .Y(_8154_)
);

AND2X2 _14392_ (
    .A(_3687_),
    .B(_3686_),
    .Y(_3672_[7])
);

FILL FILL279680x0 (
);

DFFSR _8707_ (
    .CLK(clk_bF$buf43),
    .D(_69_[25]),
    .Q(\datapath_1.regfile_1.regOut[2] [25]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL332880x286520 (
);

NAND2X1 _12705_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .B(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2270_)
);

FILL FILL68400x256880 (
);

FILL FILL272840x54340 (
);

AND2X2 _15597_ (
    .A(_4230__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_4550_)
);

AND2X2 _15177_ (
    .A(_4134_),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_4135_)
);

FILL FILL_1__8449_ (
);

FILL FILL459800x172900 (
);

FILL FILL_0__16253_ (
);

FILL FILL_1__9810_ (
);

OR2X2 _8880_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_225_)
);

OR2X2 _8460_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_5_)
);

OR2X2 _11097_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_1363_)
);

FILL FILL209760x311220 (
);

FILL FILL294880x266760 (
);

FILL FILL_0__17878_ (
);

FILL FILL_0__17458_ (
);

AND2X2 _17743_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_6663_)
);

AND2X2 _17323_ (
    .A(_6209_),
    .B(_6214_),
    .Y(_6249_)
);

FILL FILL_0__12593_ (
);

FILL FILL151240x4940 (
);

AND2X2 _9665_ (
    .A(_628_),
    .B(_627_),
    .Y(_597_[15])
);

FILL FILL129200x276640 (
);

AND2X2 _9245_ (
    .A(_408_),
    .B(_407_),
    .Y(_399_[4])
);

FILL FILL441560x88920 (
);

FILL FILL_0__8920_ (
);

FILL FILL298680x187720 (
);

FILL FILL_0__8500_ (
);

OR2X2 _18948_ (
    .A(_7849_),
    .B(_7848_),
    .Y(_7850_)
);

AND2X2 _18528_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_7436_)
);

AND2X2 _18108_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_7023_)
);

FILL FILL_1_BUFX2_insert1021 (
);

FILL FILL436240x103740 (
);

FILL FILL_1_BUFX2_insert1023 (
);

OR2X2 _13663_ (
    .A(_3146_),
    .B(_3147_),
    .Y(_3148_)
);

AND2X2 _13243_ (
    .A(_2788_),
    .B(_2780_),
    .Y(_2789_)
);

FILL FILL252320x360620 (
);

FILL FILL392920x143260 (
);

FILL FILL430160x256880 (
);

FILL FILL478800x158080 (
);

FILL FILL197600x103740 (
);

FILL FILL357960x306280 (
);

DFFSR _14868_ (
    .CLK(clk_bF$buf65),
    .D(_3870_[16]),
    .Q(_2_[16]),
    .R(rst_bF$buf26),
    .S(vdd)
);

OR2X2 _14448_ (
    .A(memoryOutData[26]),
    .B(_3737__bF$buf0),
    .Y(_3725_)
);

OR2X2 _14028_ (
    .A(_3443_),
    .B(_3442_),
    .Y(_3444_)
);

FILL FILL_1__16951_ (
);

FILL FILL191520x256880 (
);

FILL FILL_0__15524_ (
);

FILL FILL_0__15104_ (
);

FILL FILL298680x64220 (
);

AND2X2 _18281_ (
    .A(_6293__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_7193_)
);

FILL FILL64600x286520 (
);

FILL FILL387600x360620 (
);

OR2X2 _10788_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_1197_)
);

DFFSR _10368_ (
    .CLK(clk_bF$buf75),
    .D(_927_[9]),
    .Q(\datapath_1.regfile_1.regOut[15] [9]),
    .R(rst_bF$buf27),
    .S(vdd)
);

FILL FILL_0__16729_ (
);

FILL FILL_0__16309_ (
);

FILL FILL247760x345800 (
);

AND2X2 _19486_ (
    .A(_8359_),
    .B(_8358_),
    .Y(_8320_[19])
);

AND2X2 _19066_ (
    .A(_6282__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [26]),
    .Y(_7966_)
);

AND2X2 _8936_ (
    .A(_262_),
    .B(_261_),
    .Y(_201_[30])
);

AND2X2 _8516_ (
    .A(_42_),
    .B(_41_),
    .Y(_3_[19])
);

FILL FILL500840x4940 (
);

FILL FILL_1_BUFX2_insert641 (
);

OR2X2 _12934_ (
    .A(_2375_),
    .B(_2378_),
    .Y(_2498_)
);

FILL FILL_0__12649_ (
);

FILL FILL_1_BUFX2_insert643 (
);

OR2X2 _12514_ (
    .A(_2106_),
    .B(_0_),
    .Y(IorD)
);

FILL FILL_0__12229_ (
);

FILL FILL104880x360620 (
);

FILL FILL339720x281580 (
);

FILL FILL22800x148200 (
);

FILL FILL345800x222300 (
);

FILL FILL_0__16482_ (
);

FILL FILL_0__16062_ (
);

FILL FILL41040x217360 (
);

FILL FILL284240x158080 (
);

FILL FILL371640x163020 (
);

OR2X2 _13719_ (
    .A(_3194_),
    .B(_3195_),
    .Y(_3196_)
);

FILL FILL22040x375440 (
);

FILL FILL_1__15802_ (
);

FILL FILL3800x4940 (
);

FILL FILL_1__18274_ (
);

BUFX2 BUFX2_insert310 (
    .A(_68_),
    .Y(_68__bF$buf2)
);

BUFX2 BUFX2_insert311 (
    .A(_68_),
    .Y(_68__bF$buf1)
);

BUFX2 BUFX2_insert312 (
    .A(_68_),
    .Y(_68__bF$buf0)
);

BUFX2 BUFX2_insert313 (
    .A(_3869_),
    .Y(_3869__bF$buf4)
);

AND2X2 _17972_ (
    .A(_6326__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_6889_)
);

BUFX2 BUFX2_insert314 (
    .A(_3869_),
    .Y(_3869__bF$buf3)
);

BUFX2 BUFX2_insert315 (
    .A(_3869_),
    .Y(_3869__bF$buf2)
);

AND2X2 _17552_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [3]),
    .Y(_6475_)
);

BUFX2 BUFX2_insert316 (
    .A(_3869_),
    .Y(_3869__bF$buf1)
);

AND2X2 _17132_ (
    .A(_4236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_6061_)
);

BUFX2 BUFX2_insert317 (
    .A(_3869_),
    .Y(_3869__bF$buf0)
);

BUFX2 BUFX2_insert318 (
    .A(_464_),
    .Y(_464__bF$buf4)
);

BUFX2 BUFX2_insert319 (
    .A(_464_),
    .Y(_464__bF$buf3)
);

FILL FILL304760x44460 (
);

OR2X2 _9894_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_741_)
);

DFFSR _9474_ (
    .CLK(clk_bF$buf3),
    .D(_465_[18]),
    .Q(\datapath_1.regfile_1.regOut[8] [18]),
    .R(rst_bF$buf11),
    .S(vdd)
);

OR2X2 _9054_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_321_)
);

FILL FILL_0__10715_ (
);

AND2X2 _18757_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_7662_)
);

AND2X2 _18337_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_7248_)
);

FILL FILL117040x59280 (
);

OR2X2 _13892_ (
    .A(\datapath_1.a [25]),
    .B(_3342__bF$buf3),
    .Y(_3328_)
);

FILL FILL_0__13187_ (
);

OR2X2 _13472_ (
    .A(\datapath_1.PCJump [18]),
    .B(RegDst),
    .Y(_3004_)
);

FILL FILL202920x103740 (
);

AND2X2 _13052_ (
    .A(_2593_),
    .B(_2266_),
    .Y(_2609_)
);

FILL FILL_0__19413_ (
);

FILL FILL_1__12927_ (
);

FILL FILL_1__12507_ (
);

FILL FILL497800x138320 (
);

FILL FILL_0__9934_ (
);

AND2X2 _14677_ (
    .A(_3837_),
    .B(_3836_),
    .Y(_3804_[16])
);

AND2X2 _14257_ (
    .A(_3617_),
    .B(_3616_),
    .Y(_3606_[5])
);

FILL FILL_0__15753_ (
);

FILL FILL9880x365560 (
);

FILL FILL155800x4940 (
);

FILL FILL191520x9880 (
);

FILL FILL328320x59280 (
);

OR2X2 _18090_ (
    .A(_7004_),
    .B(_6991_),
    .Y(_7005_)
);

FILL FILL218880x79040 (
);

FILL FILL117800x187720 (
);

OR2X2 _10597_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_1124__bF$buf0),
    .Y(_1110_)
);

OR2X2 _10177_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .B(_926__bF$buf2),
    .Y(_890_)
);

FILL FILL_1__17125_ (
);

FILL FILL_1__12680_ (
);

FILL FILL_0__16958_ (
);

OR2X2 _16823_ (
    .A(_5756_),
    .B(_5749_),
    .Y(_5757_)
);

OR2X2 _16403_ (
    .A(_5342_),
    .B(_5341_),
    .Y(_5343_)
);

FILL FILL_0__16118_ (
);

AND2X2 _19295_ (
    .A(_8191_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd1 [29])
);

OR2X2 _8745_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_155_)
);

FILL FILL201400x44460 (
);

FILL FILL335920x177840 (
);

OR2X2 _17608_ (
    .A(_6529_),
    .B(_6528_),
    .Y(_6530_)
);

FILL FILL_0__12878_ (
);

AND2X2 _12743_ (
    .A(_2307_),
    .B(_2305_),
    .Y(_2308_)
);

FILL FILL_0__12458_ (
);

DFFSR _12323_ (
    .CLK(clk_bF$buf76),
    .D(_1917_[29]),
    .Q(\datapath_1.regfile_1.regOut[30] [29]),
    .R(rst_bF$buf110),
    .S(vdd)
);

FILL FILL222680x83980 (
);

FILL FILL367080x192660 (
);

FILL FILL371640x256880 (
);

FILL FILL446880x0 (
);

OR2X2 _13948_ (
    .A(_3373_),
    .B(_3374_),
    .Y(_3375_)
);

OR2X2 _13528_ (
    .A(IorD_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [13]),
    .Y(_3040_)
);

NAND2X1 _13108_ (
    .A(_2547_),
    .B(_2661_),
    .Y(_2662_)
);

FILL FILL111720x128440 (
);

FILL FILL394440x340860 (
);

FILL FILL_0__17496_ (
);

OR2X2 _17781_ (
    .A(_6693_),
    .B(_6700_),
    .Y(_6701_)
);

FILL FILL205200x44460 (
);

FILL FILL_0__17076_ (
);

AND2X2 _17361_ (
    .A(_6210_),
    .B(_6201_),
    .Y(_6287_)
);

FILL FILL_1__16816_ (
);

OR2X2 _9283_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_464__bF$buf0),
    .Y(_434_)
);

FILL FILL_0__10524_ (
);

AND2X2 _18986_ (
    .A(_6244__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_7887_)
);

AND2X2 _18566_ (
    .A(_6221__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_7474_)
);

AND2X2 _18146_ (
    .A(_6250__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_7060_)
);

FILL FILL447640x242060 (
);

AOI22X1 _13281_ (
    .A(_2229_),
    .B(_2504_),
    .C(_2548_),
    .D(_2431_),
    .Y(_2824_)
);

FILL FILL_0__19222_ (
);

FILL FILL278160x143260 (
);

FILL FILL502360x365560 (
);

FILL FILL_0__11729_ (
);

FILL FILL_0__9323_ (
);

FILL FILL_0__11309_ (
);

DFFSR _14486_ (
    .CLK(clk_bF$buf11),
    .D(_3672_[21]),
    .Q(\datapath_1.Data [21]),
    .R(rst_bF$buf36),
    .S(vdd)
);

FILL FILL411160x54340 (
);

AND2X2 _14066_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3476_)
);

FILL FILL_0__15982_ (
);

FILL FILL_0__15562_ (
);

FILL FILL_0__15142_ (
);

FILL FILL420280x271700 (
);

FILL FILL_1__17774_ (
);

FILL FILL_0__16767_ (
);

OR2X2 _16632_ (
    .A(_5568_),
    .B(_5553_),
    .Y(_5569_)
);

FILL FILL_0__16347_ (
);

AND2X2 _16212_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_5155_)
);

FILL FILL_0__11482_ (
);

FILL FILL373160x360620 (
);

OR2X2 _8974_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(_332__bF$buf0),
    .Y(_268_)
);

DFFSR _8554_ (
    .CLK(clk_bF$buf47),
    .D(_3_[1]),
    .Q(\datapath_1.regfile_1.regOut[1] [1]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL150480x79040 (
);

FILL FILL_1__18139_ (
);

FILL FILL347320x29640 (
);

OR2X2 _17837_ (
    .A(_6755_),
    .B(_6754_),
    .Y(_6756_)
);

OR2X2 _17417_ (
    .A(_6338_),
    .B(_6341_),
    .Y(_6342_)
);

NOR2X1 _12972_ (
    .A(_2533_),
    .B(_2531_),
    .Y(_2534_)
);

FILL FILL_0__12687_ (
);

AND2X2 _12552_ (
    .A(_2139_),
    .B(_2108_),
    .Y(_2140_)
);

OR2X2 _12132_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_1893_)
);

FILL FILL_0__18913_ (
);

OR2X2 _9759_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_671_)
);

DFFSR _9339_ (
    .CLK(clk_bF$buf93),
    .D(_399_[12]),
    .Q(\datapath_1.regfile_1.regOut[7] [12]),
    .R(rst_bF$buf41),
    .S(vdd)
);

FILL FILL386080x172900 (
);

FILL FILL325280x281580 (
);

OR2X2 _13757_ (
    .A(_3228_),
    .B(_3227_),
    .Y(_3229_)
);

AND2X2 _13337_ (
    .A(_2877_),
    .B(_2865_),
    .Y(_2878_)
);

FILL FILL_1__15420_ (
);

FILL FILL_0__14833_ (
);

FILL FILL_0__14413_ (
);

AND2X2 _17590_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_6513_)
);

AND2X2 _17170_ (
    .A(_4183__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_6098_)
);

FILL FILL_1__10399_ (
);

DFFSR _9092_ (
    .CLK(clk_bF$buf101),
    .D(_267_[23]),
    .Q(\datapath_1.regfile_1.regOut[5] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL_1__11760_ (
);

FILL FILL_0__15618_ (
);

OR2X2 _15903_ (
    .A(_4850_),
    .B(_4849_),
    .Y(_4851_)
);

FILL FILL_1__19097_ (
);

FILL FILL75240x306280 (
);

OR2X2 _18795_ (
    .A(_7695_),
    .B(_7698_),
    .Y(_7699_)
);

AND2X2 _18375_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_7286_)
);

FILL FILL379240x217360 (
);

NOR2X1 _13090_ (
    .A(_2644_),
    .B(_2466_),
    .Y(_2645_)
);

FILL FILL_0__19031_ (
);

FILL FILL12160x88920 (
);

FILL FILL475000x59280 (
);

FILL FILL_1__12125_ (
);

FILL FILL_0__9552_ (
);

OR2X2 _11823_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_1727_)
);

FILL FILL297160x123500 (
);

DFFSR _11403_ (
    .CLK(clk_bF$buf75),
    .D(_1455_[12]),
    .Q(\datapath_1.regfile_1.regOut[23] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

FILL FILL_0__11118_ (
);

FILL FILL65360x251940 (
);

OR2X2 _14295_ (
    .A(\datapath_1.ALUResult [18]),
    .B(_3671__bF$buf1),
    .Y(_3643_)
);

FILL FILL134520x49400 (
);

FILL FILL96520x237120 (
);

FILL FILL_0__15371_ (
);

FILL FILL206720x0 (
);

FILL FILL136040x326040 (
);

OR2X2 _12608_ (
    .A(_2172_),
    .B(_2171_),
    .Y(_2173_)
);

FILL FILL_0__16996_ (
);

FILL FILL_0__16576_ (
);

AND2X2 _16861_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_5794_)
);

OR2X2 _16441_ (
    .A(_5349_),
    .B(_5380_),
    .Y(_5381_)
);

AND2X2 _16021_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_4967_)
);

FILL FILL103360x187720 (
);

FILL FILL185440x83980 (
);

FILL FILL229520x74100 (
);

FILL FILL_1__9713_ (
);

AND2X2 _8783_ (
    .A(_180_),
    .B(_179_),
    .Y(_135_[22])
);

FILL FILL240160x247000 (
);

FILL FILL126160x271700 (
);

FILL FILL_1__18788_ (
);

FILL FILL_1__13083_ (
);

OR2X2 _17646_ (
    .A(_6567_),
    .B(_6566_),
    .Y(_6568_)
);

AND2X2 _17226_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_6153_)
);

INVX1 _12781_ (
    .A(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2346_)
);

OR2X2 _12361_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_2048__bF$buf2),
    .Y(_2006_)
);

FILL FILL_0__12076_ (
);

FILL FILL211280x9880 (
);

FILL FILL_0__18722_ (
);

DFFSR _9988_ (
    .CLK(clk_bF$buf88),
    .D(_729_[16]),
    .Q(\datapath_1.regfile_1.regOut[12] [16]),
    .R(rst_bF$buf95),
    .S(vdd)
);

OR2X2 _9568_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .B(_596__bF$buf4),
    .Y(_584_)
);

OR2X2 _9148_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_398__bF$buf1),
    .Y(_364_)
);

FILL FILL_1__11816_ (
);

FILL FILL457520x24700 (
);

FILL FILL_0__8403_ (
);

FILL FILL_0__10809_ (
);

FILL FILL_0_BUFX2_insert680 (
);

FILL FILL187720x355680 (
);

FILL FILL_0_BUFX2_insert682 (
);

FILL FILL_0_BUFX2_insert683 (
);

OR2X2 _13986_ (
    .A(_3407_),
    .B(_3406_),
    .Y(_3408_)
);

FILL FILL_0_BUFX2_insert684 (
);

FILL FILL344280x261820 (
);

FILL FILL_0_BUFX2_insert685 (
);

AND2X2 _13566_ (
    .A(_3065_),
    .B(_3064_),
    .Y(_1_[25])
);

NAND2X1 _13146_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2697_)
);

FILL FILL_0_BUFX2_insert686 (
);

FILL FILL189240x83980 (
);

FILL FILL_0_BUFX2_insert688 (
);

FILL FILL_0__19507_ (
);

FILL FILL_0__14642_ (
);

FILL FILL_0__14222_ (
);

FILL FILL15200x143260 (
);

FILL FILL274360x266760 (
);

FILL FILL434720x98800 (
);

FILL FILL488680x4940 (
);

FILL FILL_0__15847_ (
);

FILL FILL498560x103740 (
);

FILL FILL_0__15427_ (
);

OR2X2 _15712_ (
    .A(_4662_),
    .B(_4659_),
    .Y(_4663_)
);

FILL FILL_0__10982_ (
);

FILL FILL_0__10562_ (
);

OR2X2 _18184_ (
    .A(_7097_),
    .B(_7096_),
    .Y(_7098_)
);

FILL FILL145920x217360 (
);

FILL FILL492480x256880 (
);

FILL FILL_0__19260_ (
);

FILL FILL_1__17639_ (
);

FILL FILL_1__17219_ (
);

AND2X2 _16917_ (
    .A(_4172__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_5849_)
);

FILL FILL_0__9781_ (
);

FILL FILL_0__11767_ (
);

FILL FILL_0__9361_ (
);

OR2X2 _11632_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .B(_1652__bF$buf4),
    .Y(_1640_)
);

FILL FILL_0__11347_ (
);

OR2X2 _11212_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .B(_1454__bF$buf1),
    .Y(_1420_)
);

FILL FILL414200x271700 (
);

OR2X2 _19389_ (
    .A(_8276_),
    .B(_8283_),
    .Y(_8284_)
);

FILL FILL263720x88920 (
);

DFFSR _8839_ (
    .CLK(clk_bF$buf25),
    .D(_135_[28]),
    .Q(\datapath_1.regfile_1.regOut[3] [28]),
    .R(rst_bF$buf55),
    .S(vdd)
);

BUFX2 _8419_ (
    .A(_1_[27]),
    .Y(memoryAddress[27])
);

FILL FILL_0__15180_ (
);

FILL FILL_1__13979_ (
);

XOR2X1 _12837_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2402_)
);

FILL FILL266760x281580 (
);

OR2X2 _12417_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_2043_)
);

FILL FILL272840x222300 (
);

FILL FILL72200x340860 (
);

FILL FILL_0__13913_ (
);

FILL FILL_1__17392_ (
);

AND2X2 _16670_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_5606_)
);

AND2X2 _16250_ (
    .A(_5192_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd2 [15])
);

FILL FILL8360x301340 (
);

OR2X2 _8592_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_73_)
);

FILL FILL_1__10840_ (
);

FILL FILL67640x138320 (
);

FILL FILL494000x148200 (
);

FILL FILL207480x133380 (
);

AND2X2 _17875_ (
    .A(_6317__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_6793_)
);

OR2X2 _17455_ (
    .A(_6379_),
    .B(_6376_),
    .Y(_6380_)
);

FILL FILL270560x296400 (
);

AND2X2 _17035_ (
    .A(_4172__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_5965_)
);

INVX1 _12590_ (
    .A(gnd),
    .Y(_2155_)
);

DFFSR _12170_ (
    .CLK(clk_bF$buf14),
    .D(_1851_[5]),
    .Q(\datapath_1.regfile_1.regOut[29] [5]),
    .R(rst_bF$buf8),
    .S(vdd)
);

FILL FILL_0__18531_ (
);

FILL FILL_0__18111_ (
);

FILL FILL445360x335920 (
);

AND2X2 _9797_ (
    .A(_696_),
    .B(_695_),
    .Y(_663_[16])
);

AND2X2 _9377_ (
    .A(_476_),
    .B(_475_),
    .Y(_465_[5])
);

FILL FILL_1__11205_ (
);

FILL FILL133000x360620 (
);

FILL FILL_0__8632_ (
);

DFFSR _10903_ (
    .CLK(clk_bF$buf84),
    .D(_1191_[28]),
    .Q(\datapath_1.regfile_1.regOut[19] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL351120x163020 (
);

AND2X2 _13795_ (
    .A(_3084__bF$buf4),
    .B(\datapath_1.PCJump [29]),
    .Y(_3261_)
);

NAND3X1 _13375_ (
    .A(_2383_),
    .B(_2912_),
    .C(_2908_),
    .Y(_2913_)
);

FILL FILL388360x286520 (
);

FILL FILL160360x316160 (
);

FILL FILL302480x350740 (
);

FILL FILL_0__9837_ (
);

FILL FILL289560x98800 (
);

FILL FILL482600x242060 (
);

FILL FILL_1__16243_ (
);

FILL FILL437000x365560 (
);

FILL FILL215840x9880 (
);

AND2X2 _15941_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_4888_)
);

AND2X2 _15521_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_4475_)
);

FILL FILL_0__15236_ (
);

AND2X2 _15101_ (
    .A(_4074_),
    .B(_4083_),
    .Y(\datapath_1.regfile_1.regEn [7])
);

FILL FILL_0__10791_ (
);

FILL FILL385320x182780 (
);

FILL FILL_1__17868_ (
);

FILL FILL234840x9880 (
);

OR2X2 _16726_ (
    .A(_5659_),
    .B(_5660_),
    .Y(_5661_)
);

OR2X2 _16306_ (
    .A(_5247_),
    .B(_5246_),
    .Y(_5248_)
);

FILL FILL332880x172900 (
);

FILL FILL_0__9170_ (
);

FILL FILL_0__11576_ (
);

AND2X2 _11861_ (
    .A(_1752_),
    .B(_1751_),
    .Y(_1719_[16])
);

AND2X2 _11441_ (
    .A(_1532_),
    .B(_1531_),
    .Y(_1521_[5])
);

DFFSR _11021_ (
    .CLK(clk_bF$buf11),
    .D(_1257_[17]),
    .Q(\datapath_1.regfile_1.regOut[20] [17]),
    .R(rst_bF$buf111),
    .S(vdd)
);

OR2X2 _19198_ (
    .A(_8094_),
    .B(_8095_),
    .Y(_8096_)
);

FILL FILL281960x340860 (
);

FILL FILL_0__17802_ (
);

AND2X2 _8648_ (
    .A(_110_),
    .B(_109_),
    .Y(_69_[20])
);

FILL FILL_1__13368_ (
);

XNOR2X1 _12646_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2211_)
);

OR2X2 _12226_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .B(_1982__bF$buf0),
    .Y(_1936_)
);

FILL FILL_0__13722_ (
);

FILL FILL_0_BUFX2_insert1031 (
);

FILL FILL_0_BUFX2_insert1033 (
);

FILL FILL_0__16194_ (
);

FILL FILL_0_BUFX2_insert1035 (
);

FILL FILL_0_BUFX2_insert1037 (
);

FILL FILL_0_BUFX2_insert1038 (
);

FILL FILL_0_BUFX2_insert1039 (
);

FILL FILL99560x340860 (
);

FILL FILL334400x340860 (
);

FILL FILL370120x98800 (
);

FILL FILL_0__14927_ (
);

FILL FILL_0__17399_ (
);

OR2X2 _17684_ (
    .A(_6604_),
    .B(_6603_),
    .Y(_6605_)
);

AND2X2 _17264_ (
    .A(_4183__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_6191_)
);

FILL FILL_0__18760_ (
);

FILL FILL_0__18340_ (
);

FILL FILL277400x291460 (
);

OR2X2 _9186_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_389_)
);

FILL FILL374680x242060 (
);

FILL FILL_0__8861_ (
);

FILL FILL_0__10847_ (
);

FILL FILL_0__8441_ (
);

AND2X2 _10712_ (
    .A(_1166_),
    .B(_1165_),
    .Y(_1125_[20])
);

FILL FILL_0__10427_ (
);

FILL FILL_0__10007_ (
);

OR2X2 _18889_ (
    .A(_7791_),
    .B(_7789_),
    .Y(_7792_)
);

NOR2X1 _18469_ (
    .A(_6310__bF$buf4),
    .B(_7377_),
    .Y(_7378_)
);

AND2X2 _18049_ (
    .A(_6250__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_6965_)
);

OR2X2 _13184_ (
    .A(_2418_),
    .B(_2732_),
    .Y(_2733_)
);

FILL FILL181640x59280 (
);

AND2X2 _19410_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_8305_)
);

FILL FILL_0__19125_ (
);

FILL FILL_0__14680_ (
);

FILL FILL_1__12219_ (
);

FILL FILL_0__9646_ (
);

DFFSR _11917_ (
    .CLK(clk_bF$buf33),
    .D(_1719_[10]),
    .Q(\datapath_1.regfile_1.regOut[27] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

AND2X2 _14389_ (
    .A(_3685_),
    .B(_3684_),
    .Y(_3672_[6])
);

FILL FILL_1__16892_ (
);

FILL FILL123120x103740 (
);

FILL FILL_1__16472_ (
);

AND2X2 _15750_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_4700_)
);

FILL FILL_0__15465_ (
);

FILL FILL_0__15045_ (
);

AND2X2 _15330_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_4287_)
);

FILL FILL_1__17257_ (
);

FILL FILL395960x360620 (
);

AND2X2 _16955_ (
    .A(_4234__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_5886_)
);

OR2X2 _16535_ (
    .A(_5469_),
    .B(_5472_),
    .Y(_5473_)
);

AND2X2 _16115_ (
    .A(_4241__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_5060_)
);

DFFSR _11670_ (
    .CLK(clk_bF$buf43),
    .D(_1587_[21]),
    .Q(\datapath_1.regfile_1.regOut[25] [21]),
    .R(rst_bF$buf41),
    .S(vdd)
);

OR2X2 _11250_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_1445_)
);

FILL FILL_0__17611_ (
);

FILL FILL427120x108680 (
);

OR2X2 _8877_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_223_)
);

INVX2 _8457_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .Y(_68_)
);

FILL FILL_1__13597_ (
);

FILL FILL129200x39520 (
);

FILL FILL5320x158080 (
);

OR2X2 _12875_ (
    .A(_2439_),
    .B(_2422_),
    .Y(_2440_)
);

FILL FILL_1__19403_ (
);

INVX1 _12455_ (
    .A(\aluControl_1.inst [3]),
    .Y(_2049_)
);

AND2X2 _12035_ (
    .A(_1848_),
    .B(_1847_),
    .Y(_1785_[31])
);

FILL FILL_0__13531_ (
);

FILL FILL_0__13111_ (
);

FILL FILL481080x34580 (
);

FILL FILL_0__8917_ (
);

FILL FILL_1__9560_ (
);

FILL FILL_0__14316_ (
);

DFFSR _14601_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[7]),
    .Q(\datapath_1.PCJump [9]),
    .R(rst_bF$buf100),
    .S(vdd)
);

FILL FILL160360x39520 (
);

AND2X2 _17493_ (
    .A(_6206__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_6417_)
);

AND2X2 _17073_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_6003_)
);

FILL FILL123880x232180 (
);

FILL FILL335160x49400 (
);

FILL FILL_1__16108_ (
);

AND2X2 _15806_ (
    .A(_4197__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_4755_)
);

FILL FILL15200x306280 (
);

FILL FILL_0__8670_ (
);

OR2X2 _10941_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_1279_)
);

FILL FILL_0__10656_ (
);

INVX2 _10521_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .Y(_1124_)
);

DFFSR _10101_ (
    .CLK(clk_bF$buf96),
    .D(_795_[0]),
    .Q(\datapath_1.regfile_1.regOut[13] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL8360x54340 (
);

OR2X2 _18698_ (
    .A(_7603_),
    .B(_7600_),
    .Y(_7604_)
);

OR2X2 _18278_ (
    .A(_7189_),
    .B(_7188_),
    .Y(_7190_)
);

FILL FILL_0__19354_ (
);

FILL FILL_0__9875_ (
);

FILL FILL_0__9455_ (
);

FILL FILL_0__9035_ (
);

AND2X2 _11726_ (
    .A(_1682_),
    .B(_1681_),
    .Y(_1653_[14])
);

FILL FILL164160x39520 (
);

AND2X2 _11306_ (
    .A(_1462_),
    .B(_1461_),
    .Y(_1455_[3])
);

FILL FILL442320x301340 (
);

OR2X2 _14198_ (
    .A(\datapath_1.Data [18]),
    .B(_3605__bF$buf4),
    .Y(_3577_)
);

FILL FILL291840x54340 (
);

FILL FILL_0__15694_ (
);

FILL FILL372400x306280 (
);

FILL FILL313880x355680 (
);

FILL FILL13680x365560 (
);

FILL FILL_0__16479_ (
);

AND2X2 _16764_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_5698_)
);

FILL FILL_0__16059_ (
);

OR2X2 _16344_ (
    .A(_5277_),
    .B(_5284_),
    .Y(_5285_)
);

FILL FILL_0__17840_ (
);

FILL FILL_0__17000_ (
);

DFFSR _8686_ (
    .CLK(clk_bF$buf87),
    .D(_69_[4]),
    .Q(\datapath_1.regfile_1.regOut[2] [4]),
    .R(rst_bF$buf2),
    .S(vdd)
);

BUFX2 BUFX2_insert280 (
    .A(_3605_),
    .Y(_3605__bF$buf2)
);

BUFX2 BUFX2_insert281 (
    .A(_3605_),
    .Y(_3605__bF$buf1)
);

BUFX2 BUFX2_insert282 (
    .A(_3605_),
    .Y(_3605__bF$buf0)
);

BUFX2 BUFX2_insert283 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf4 )
);

BUFX2 BUFX2_insert284 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf3 )
);

AND2X2 _17969_ (
    .A(_6297__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_6886_)
);

BUFX2 BUFX2_insert285 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf2 )
);

AND2X2 _17549_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_6472_)
);

BUFX2 BUFX2_insert286 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf1 )
);

AND2X2 _17129_ (
    .A(_4200__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_6058_)
);

BUFX2 BUFX2_insert287 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf0 )
);

BUFX2 BUFX2_insert288 (
    .A(_4181_),
    .Y(_4181__bF$buf4)
);

OR2X2 _12684_ (
    .A(_2246_),
    .B(_2248_),
    .Y(_2249_)
);

BUFX2 BUFX2_insert289 (
    .A(_4181_),
    .Y(_4181__bF$buf3)
);

OR2X2 _12264_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_1961_)
);

FILL FILL86640x24700 (
);

FILL FILL_0__18625_ (
);

AND2X2 _18910_ (
    .A(_6315__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_7812_)
);

FILL FILL_0__18205_ (
);

FILL FILL_0__13760_ (
);

FILL FILL_0__13340_ (
);

FILL FILL279680x256880 (
);

FILL FILL_0__8726_ (
);

FILL FILL85880x113620 (
);

OR2X2 _13889_ (
    .A(\datapath_1.a [24]),
    .B(_3342__bF$buf0),
    .Y(_3326_)
);

AND2X2 _13469_ (
    .A(_3001_),
    .B(_2561_),
    .Y(_3002_)
);

XNOR2X1 _13049_ (
    .A(_2267_),
    .B(_2605_),
    .Y(_2606_)
);

FILL FILL66880x271700 (
);

FILL FILL_0__14965_ (
);

AND2X2 _14830_ (
    .A(_3919_),
    .B(_3918_),
    .Y(_3870_[24])
);

FILL FILL_0__14545_ (
);

AND2X2 _14410_ (
    .A(_3699_),
    .B(_3698_),
    .Y(_3672_[13])
);

FILL FILL231800x276640 (
);

FILL FILL_1__16757_ (
);

FILL FILL_1__16337_ (
);

FILL FILL_1__11892_ (
);

AND2X2 _15615_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_4567_)
);

DFFSR _10750_ (
    .CLK(clk_bF$buf82),
    .D(_1125_[4]),
    .Q(\datapath_1.regfile_1.regOut[18] [4]),
    .R(rst_bF$buf94),
    .S(vdd)
);

FILL FILL_0__10045_ (
);

OR2X2 _10330_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .B(_992__bF$buf0),
    .Y(_972_)
);

OR2X2 _18087_ (
    .A(_7001_),
    .B(_7000_),
    .Y(_7002_)
);

FILL FILL_0__19163_ (
);

FILL FILL_1__12257_ (
);

FILL FILL_0__9684_ (
);

OR2X2 _11955_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_1795_)
);

DFFSR _11535_ (
    .CLK(clk_bF$buf48),
    .D(_1521_[15]),
    .Q(\datapath_1.regfile_1.regOut[24] [15]),
    .R(rst_bF$buf21),
    .S(vdd)
);

OR2X2 _11115_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_1375_)
);

FILL FILL193800x256880 (
);

FILL FILL_0__12611_ (
);

FILL FILL_0__15083_ (
);

FILL FILL_1__8640_ (
);

FILL FILL212800x222300 (
);

FILL FILL_1__14403_ (
);

FILL FILL_0__13816_ (
);

FILL FILL151240x158080 (
);

AND2X2 _16993_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_5924_)
);

OR2X2 _16573_ (
    .A(_5508_),
    .B(_5509_),
    .Y(_5510_)
);

FILL FILL_0__16288_ (
);

OR2X2 _16153_ (
    .A(_5096_),
    .B(_5081_),
    .Y(_5097_)
);

FILL FILL_1__9005_ (
);

FILL FILL413440x202540 (
);

AND2X2 _8495_ (
    .A(_28_),
    .B(_27_),
    .Y(_3_[12])
);

FILL FILL298680x370500 (
);

AND2X2 _17778_ (
    .A(_6264__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_6698_)
);

AND2X2 _17358_ (
    .A(_6272__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_6284_)
);

FILL FILL210520x296400 (
);

AND2X2 _12493_ (
    .A(_2091_),
    .B(\control_1.reg_state.dout [1]),
    .Y(_2096_)
);

OR2X2 _12073_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .B(_1916__bF$buf4),
    .Y(_1854_)
);

FILL FILL_1__19021_ (
);

FILL FILL207480x247000 (
);

FILL FILL_0__18854_ (
);

FILL FILL43320x217360 (
);

FILL FILL430160x118560 (
);

FILL FILL_1__11948_ (
);

FILL FILL56240x163020 (
);

OR2X2 _10806_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_1209_)
);

FILL FILL367840x0 (
);

FILL FILL60800x227240 (
);

OR2X2 _13698_ (
    .A(_3176_),
    .B(_3177_),
    .Y(_3178_)
);

AND2X2 _13278_ (
    .A(_2820_),
    .B(_2423_),
    .Y(_2821_)
);

FILL FILL_1__15361_ (
);

FILL FILL_0__19219_ (
);

AND2X2 _19504_ (
    .A(_8371_),
    .B(_8370_),
    .Y(_8320_[25])
);

FILL FILL_0__14774_ (
);

FILL FILL451440x370500 (
);

FILL FILL_1__16986_ (
);

FILL FILL_0__15979_ (
);

AND2X2 _15844_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_4793_)
);

FILL FILL_0__15559_ (
);

OR2X2 _15424_ (
    .A(_4377_),
    .B(_4378_),
    .Y(_4379_)
);

DFFSR _15004_ (
    .CLK(clk_bF$buf77),
    .D(_3936_[23]),
    .Q(\datapath_1.mux_iord.din0 [23]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL104120x237120 (
);

FILL FILL_0__16920_ (
);

FILL FILL_0__16500_ (
);

FILL FILL156560x34580 (
);

FILL FILL235600x316160 (
);

OR2X2 _16629_ (
    .A(_5565_),
    .B(_5564_),
    .Y(_5566_)
);

AND2X2 _16209_ (
    .A(_4214__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_5152_)
);

FILL FILL_0__9493_ (
);

FILL FILL_0__11899_ (
);

FILL FILL_0__11479_ (
);

OR2X2 _11764_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .B(_1718__bF$buf4),
    .Y(_1708_)
);

FILL FILL_0__11059_ (
);

OR2X2 _11344_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .B(_1520__bF$buf3),
    .Y(_1488_)
);

FILL FILL465880x29640 (
);

FILL FILL_0__17705_ (
);

FILL FILL_0__12840_ (
);

FILL FILL_0__12420_ (
);

OR2X2 _9912_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_753_)
);

MUX2X1 _12969_ (
    .A(_2501_),
    .B(_2376__bF$buf3),
    .S(_2358_),
    .Y(_2531_)
);

OR2X2 _12549_ (
    .A(_2131_),
    .B(_2137_),
    .Y(\control_1.next [1])
);

OR2X2 _12129_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_1891_)
);

FILL FILL_1_BUFX2_insert995 (
);

FILL FILL_1_BUFX2_insert997 (
);

FILL FILL_1__14212_ (
);

FILL FILL_1_BUFX2_insert999 (
);

OR2X2 _13910_ (
    .A(\datapath_1.a [31]),
    .B(_3342__bF$buf4),
    .Y(_3340_)
);

FILL FILL_0__13205_ (
);

FILL FILL362520x321100 (
);

AND2X2 _16382_ (
    .A(_4158__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_5322_)
);

FILL FILL114760x64220 (
);

FILL FILL_1__15837_ (
);

FILL FILL_1__10972_ (
);

BUFX2 BUFX2_insert660 (
    .A(_6300_),
    .Y(_6300__bF$buf4)
);

BUFX2 BUFX2_insert661 (
    .A(_6300_),
    .Y(_6300__bF$buf3)
);

BUFX2 BUFX2_insert662 (
    .A(_6300_),
    .Y(_6300__bF$buf2)
);

BUFX2 BUFX2_insert663 (
    .A(_6300_),
    .Y(_6300__bF$buf1)
);

FILL FILL133000x19760 (
);

BUFX2 BUFX2_insert664 (
    .A(_6300_),
    .Y(_6300__bF$buf0)
);

AND2X2 _17587_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_6510_)
);

BUFX2 BUFX2_insert665 (
    .A(_860_),
    .Y(_860__bF$buf4)
);

BUFX2 BUFX2_insert666 (
    .A(_860_),
    .Y(_860__bF$buf3)
);

OR2X2 _17167_ (
    .A(_6094_),
    .B(_6093_),
    .Y(_6095_)
);

BUFX2 BUFX2_insert667 (
    .A(_860_),
    .Y(_860__bF$buf2)
);

BUFX2 BUFX2_insert668 (
    .A(_860_),
    .Y(_860__bF$buf1)
);

BUFX2 BUFX2_insert669 (
    .A(_860_),
    .Y(_860__bF$buf0)
);

FILL FILL369360x192660 (
);

FILL FILL78280x0 (
);

FILL FILL_0__18243_ (
);

DFFSR _9089_ (
    .CLK(clk_bF$buf9),
    .D(_267_[20]),
    .Q(\datapath_1.regfile_1.regOut[5] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

FILL FILL389880x44460 (
);

FILL FILL_1__11337_ (
);

FILL FILL75240x34580 (
);

FILL FILL_0__8764_ (
);

OR2X2 _10615_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .B(_1124__bF$buf4),
    .Y(_1122_)
);

FILL FILL396720x340860 (
);

NAND2X1 _13087_ (
    .A(_2641_),
    .B(_2640_),
    .Y(_2642_)
);

FILL FILL_1__15590_ (
);

FILL FILL_0__19448_ (
);

FILL FILL_0__19028_ (
);

AND2X2 _19313_ (
    .A(_6247__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_8209_)
);

FILL FILL228000x44460 (
);

FILL FILL_0__14163_ (
);

FILL FILL19000x14820 (
);

FILL FILL_0__9969_ (
);

FILL FILL_0__9129_ (
);

FILL FILL_1__13903_ (
);

FILL FILL_0__15788_ (
);

AND2X2 _15653_ (
    .A(_4130__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_4605_)
);

OR2X2 _15233_ (
    .A(_4190_),
    .B(_4188_),
    .Y(_4191_)
);

FILL FILL174800x69160 (
);

FILL FILL504640x365560 (
);

FILL FILL248520x355680 (
);

FILL FILL18240x360620 (
);

AND2X2 _16858_ (
    .A(_4181__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [25]),
    .Y(_5791_)
);

OR2X2 _16438_ (
    .A(_5374_),
    .B(_5377_),
    .Y(_5378_)
);

FILL FILL354160x108680 (
);

AND2X2 _16018_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_4964_)
);

AND2X2 _11993_ (
    .A(_1820_),
    .B(_1819_),
    .Y(_1785_[17])
);

FILL FILL_1__18521_ (
);

AND2X2 _11573_ (
    .A(_1600_),
    .B(_1599_),
    .Y(_1587_[6])
);

FILL FILL_1__18101_ (
);

DFFSR _11153_ (
    .CLK(clk_bF$buf46),
    .D(_1323_[20]),
    .Q(\datapath_1.regfile_1.regOut[21] [20]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _9721_ (
    .CLK(clk_bF$buf29),
    .D(_597_[7]),
    .Q(\datapath_1.regfile_1.regOut[10] [7]),
    .R(rst_bF$buf21),
    .S(vdd)
);

OR2X2 _9301_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .B(_464__bF$buf4),
    .Y(_446_)
);

OR2X2 _12778_ (
    .A(_2326_),
    .B(_2342_),
    .Y(_2343_)
);

OR2X2 _12358_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_2048__bF$buf4),
    .Y(_2004_)
);

FILL FILL_0__18719_ (
);

FILL FILL_0__13854_ (
);

FILL FILL_0__13434_ (
);

AND2X2 _16191_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_5134_)
);

FILL FILL37240x64220 (
);

FILL FILL_1__15226_ (
);

OR2X2 _14924_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [13]),
    .Y(_3962_)
);

FILL FILL_0__14219_ (
);

OR2X2 _14504_ (
    .A(IRWrite_bF$buf4),
    .B(\aluControl_1.inst [2]),
    .Y(_3742_)
);

FILL FILL12160x301340 (
);

AND2X2 _17396_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_6322_)
);

FILL FILL388360x172900 (
);

FILL FILL316160x212420 (
);

FILL FILL_0__18892_ (
);

FILL FILL_0__18472_ (
);

FILL FILL_0__18052_ (
);

FILL FILL327560x281580 (
);

AND2X2 _15709_ (
    .A(_4142__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_4660_)
);

FILL FILL_0__8993_ (
);

AND2X2 _10844_ (
    .A(_1234_),
    .B(_1233_),
    .Y(_1191_[21])
);

FILL FILL_0__10559_ (
);

FILL FILL_0__10139_ (
);

AND2X2 _10424_ (
    .A(_1014_),
    .B(_1013_),
    .Y(_993_[10])
);

OR2X2 _10004_ (
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .Y(_859_)
);

FILL FILL_0__11500_ (
);

DFFSR _19542_ (
    .CLK(clk_bF$buf80),
    .D(_8320_[19]),
    .Q(\datapath_1.regfile_1.regOut[0] [19]),
    .R(rst_bF$buf76),
    .S(vdd)
);

AND2X2 _19122_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_8021_)
);

FILL FILL95000x133380 (
);

FILL FILL418000x24700 (
);

FILL FILL164160x123500 (
);

FILL FILL132240x335920 (
);

FILL FILL_0__9778_ (
);

OR2X2 _11629_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .B(_1652__bF$buf0),
    .Y(_1638_)
);

OR2X2 _11209_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .B(_1454__bF$buf2),
    .Y(_1418_)
);

FILL FILL_0__12705_ (
);

FILL FILL58520x88920 (
);

FILL FILL_0__15597_ (
);

AND2X2 _15882_ (
    .A(_4158__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_4830_)
);

OR2X2 _15462_ (
    .A(_4416_),
    .B(_4415_),
    .Y(_4417_)
);

FILL FILL_0__15177_ (
);

INVX1 _15042_ (
    .A(_4003_),
    .Y(_4031_)
);

FILL FILL202920x59280 (
);

AND2X2 _16667_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_5603_)
);

OR2X2 _16247_ (
    .A(_5182_),
    .B(_5189_),
    .Y(_5190_)
);

FILL FILL_1__18750_ (
);

FILL FILL120840x108680 (
);

OR2X2 _11382_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_1513_)
);

FILL FILL_0__17743_ (
);

FILL FILL_0__17323_ (
);

FILL FILL221160x316160 (
);

OR2X2 _8589_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_71_)
);

FILL FILL228000x192660 (
);

AND2X2 _9950_ (
    .A(_778_),
    .B(_777_),
    .Y(_729_[24])
);

AND2X2 _9530_ (
    .A(_558_),
    .B(_557_),
    .Y(_531_[13])
);

AND2X2 _9110_ (
    .A(_338_),
    .B(_337_),
    .Y(_333_[2])
);

DFFSR _12587_ (
    .CLK(clk_bF$buf20),
    .D(_2143_[3]),
    .Q(\control_1.reg_state.dout [3]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _12167_ (
    .CLK(clk_bF$buf112),
    .D(_1851_[2]),
    .Q(\datapath_1.regfile_1.regOut[29] [2]),
    .R(rst_bF$buf3),
    .S(vdd)
);

FILL FILL_1__14250_ (
);

FILL FILL_0__18948_ (
);

OR2X2 _18813_ (
    .A(_7716_),
    .B(_7713_),
    .Y(_7717_)
);

FILL FILL_0_BUFX2_insert300 (
);

FILL FILL_0__18108_ (
);

FILL FILL_0_BUFX2_insert302 (
);

FILL FILL_0_BUFX2_insert303 (
);

FILL FILL_0_BUFX2_insert304 (
);

FILL FILL_0_BUFX2_insert305 (
);

FILL FILL_0_BUFX2_insert306 (
);

FILL FILL_0_BUFX2_insert307 (
);

FILL FILL_0_BUFX2_insert309 (
);

FILL FILL269040x24700 (
);

FILL FILL_1__9692_ (
);

FILL FILL242440x247000 (
);

FILL FILL452200x123500 (
);

FILL FILL_1__15875_ (
);

FILL FILL_1__15455_ (
);

FILL FILL_1__10590_ (
);

DFFSR _14733_ (
    .CLK(clk_bF$buf15),
    .D(_3804_[10]),
    .Q(\datapath_1.a [10]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL_0__14448_ (
);

FILL FILL_0__14028_ (
);

OR2X2 _14313_ (
    .A(\datapath_1.ALUResult [24]),
    .B(_3671__bF$buf3),
    .Y(_3655_)
);

FILL FILL463600x192660 (
);

FILL FILL91200x163020 (
);

FILL FILL288800x64220 (
);

FILL FILL502360x34580 (
);

FILL FILL_0__18281_ (
);

FILL FILL430160x98800 (
);

FILL FILL412680x69160 (
);

AND2X2 _15938_ (
    .A(_4181__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_4885_)
);

FILL FILL259160x256880 (
);

AND2X2 _15518_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_4472_)
);

OR2X2 _10653_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_1127_)
);

DFFSR _10233_ (
    .CLK(clk_bF$buf79),
    .D(_861_[3]),
    .Q(\datapath_1.regfile_1.regOut[14] [3]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL_0__19066_ (
);

OR2X2 _19351_ (
    .A(_8245_),
    .B(_8246_),
    .Y(_8247_)
);

FILL FILL46360x271700 (
);

AND2X2 _8801_ (
    .A(_192_),
    .B(_191_),
    .Y(_135_[28])
);

AND2X2 _11858_ (
    .A(_1750_),
    .B(_1749_),
    .Y(_1719_[15])
);

AND2X2 _11438_ (
    .A(_1530_),
    .B(_1529_),
    .Y(_1521_[4])
);

DFFSR _11018_ (
    .CLK(clk_bF$buf98),
    .D(_1257_[14]),
    .Q(\datapath_1.regfile_1.regOut[20] [14]),
    .R(rst_bF$buf87),
    .S(vdd)
);

FILL FILL_0__12934_ (
);

AND2X2 _15691_ (
    .A(_4146__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [7]),
    .Y(_4642_)
);

AND2X2 _15271_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_4229_)
);

FILL FILL_1__8543_ (
);

FILL FILL416480x69160 (
);

FILL FILL338200x291460 (
);

FILL FILL66880x4940 (
);

FILL FILL_1__17198_ (
);

OR2X2 _16896_ (
    .A(_5826_),
    .B(_5827_),
    .Y(_5828_)
);

OR2X2 _16476_ (
    .A(_5413_),
    .B(_5414_),
    .Y(_5415_)
);

OR2X2 _16056_ (
    .A(_5001_),
    .B(_4986_),
    .Y(_5002_)
);

FILL FILL340480x202540 (
);

FILL FILL380000x311220 (
);

OR2X2 _11191_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_1454__bF$buf2),
    .Y(_1406_)
);

FILL FILL452960x59280 (
);

FILL FILL_0__17972_ (
);

BUFX2 _8398_ (
    .A(_1_[6]),
    .Y(memoryAddress[6])
);

FILL FILL_1__10226_ (
);

FILL FILL38000x167960 (
);

OR2X2 _12396_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_2029_)
);

FILL FILL_0__18757_ (
);

AND2X2 _18622_ (
    .A(_6238__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_7529_)
);

FILL FILL_0__18337_ (
);

AND2X2 _18202_ (
    .A(_6297__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_7115_)
);

FILL FILL_0__13472_ (
);

FILL FILL_0__13052_ (
);

FILL FILL475760x202540 (
);

FILL FILL_0__8438_ (
);

AND2X2 _10709_ (
    .A(_1164_),
    .B(_1163_),
    .Y(_1125_[19])
);

FILL FILL316920x54340 (
);

AND2X2 _19407_ (
    .A(_6287__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_8302_)
);

AND2X2 _14962_ (
    .A(_3987_),
    .B(_3986_),
    .Y(_3936_[25])
);

FILL FILL_0__14677_ (
);

FILL FILL_0__14257_ (
);

AND2X2 _14542_ (
    .A(_3767_),
    .B(_3766_),
    .Y(_3738_[14])
);

AND2X2 _14122_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3524_)
);

FILL FILL395200x167960 (
);

FILL FILL482600x172900 (
);

FILL FILL109440x54340 (
);

FILL FILL479560x123500 (
);

FILL FILL23560x83980 (
);

FILL FILL215080x301340 (
);

FILL FILL_0__18090_ (
);

FILL FILL180120x143260 (
);

FILL FILL505400x118560 (
);

FILL FILL353400x163020 (
);

AND2X2 _15747_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_4697_)
);

OR2X2 _15327_ (
    .A(_4283_),
    .B(_4282_),
    .Y(_4284_)
);

FILL FILL_0__10597_ (
);

DFFSR _10882_ (
    .CLK(clk_bF$buf90),
    .D(_1191_[7]),
    .Q(\datapath_1.regfile_1.regOut[19] [7]),
    .R(rst_bF$buf108),
    .S(vdd)
);

OR2X2 _10462_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_1058__bF$buf1),
    .Y(_1040_)
);

FILL FILL_0__10177_ (
);

OR2X2 _10042_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .B(_860__bF$buf2),
    .Y(_820_)
);

FILL FILL_0__16823_ (
);

FILL FILL162640x316160 (
);

FILL FILL_0__19295_ (
);

FILL FILL304760x350740 (
);

OR2X2 _19160_ (
    .A(_8055_),
    .B(_8058_),
    .Y(_8059_)
);

FILL FILL477280x197600 (
);

OR2X2 _8610_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_85_)
);

FILL FILL_1__12389_ (
);

DFFSR _11667_ (
    .CLK(clk_bF$buf3),
    .D(_1587_[18]),
    .Q(\datapath_1.regfile_1.regOut[25] [18]),
    .R(rst_bF$buf58),
    .S(vdd)
);

FILL FILL_1__18615_ (
);

OR2X2 _11247_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_1443_)
);

FILL FILL142120x59280 (
);

FILL FILL_1__13330_ (
);

FILL FILL_0__17608_ (
);

FILL FILL431680x39520 (
);

NOR2X1 _15080_ (
    .A(_4049_),
    .B(_4065__bF$buf2),
    .Y(_4066_)
);

FILL FILL367840x311220 (
);

AND2X2 _9815_ (
    .A(_708_),
    .B(_707_),
    .Y(_663_[22])
);

FILL FILL_1__14535_ (
);

FILL FILL462840x9880 (
);

FILL FILL454480x222300 (
);

FILL FILL_0__13948_ (
);

OR2X2 _13813_ (
    .A(_3276_),
    .B(_3275_),
    .Y(_3277_)
);

FILL FILL_0__13528_ (
);

AND2X2 _16285_ (
    .A(_4158__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_5227_)
);

FILL FILL_0__17361_ (
);

FILL FILL133000x222300 (
);

FILL FILL481840x9880 (
);

FILL FILL_1__10035_ (
);

FILL FILL391400x197600 (
);

FILL FILL104880x182780 (
);

FILL FILL270560x345800 (
);

FILL FILL180880x44460 (
);

FILL FILL_0__18986_ (
);

FILL FILL_0__18566_ (
);

AND2X2 _18851_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_7754_)
);

FILL FILL_0__18146_ (
);

OR2X2 _18431_ (
    .A(_7332_),
    .B(_7340_),
    .Y(_7341_)
);

AND2X2 _18011_ (
    .A(_6244__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_6927_)
);

FILL FILL64600x44460 (
);

FILL FILL_0__13281_ (
);

FILL FILL19760x242060 (
);

FILL FILL465120x34580 (
);

FILL FILL355680x54340 (
);

FILL FILL_0__8667_ (
);

OR2X2 _10938_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_1277_)
);

DFFSR _10518_ (
    .CLK(clk_bF$buf108),
    .D(_993_[30]),
    .Q(\datapath_1.regfile_1.regOut[16] [30]),
    .R(rst_bF$buf93),
    .S(vdd)
);

FILL FILL351120x212420 (
);

FILL FILL86640x9880 (
);

FILL FILL124640x24700 (
);

AND2X2 _19216_ (
    .A(_6297__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_8114_)
);

OR2X2 _14771_ (
    .A(vdd),
    .B(_2_[5]),
    .Y(_3880_)
);

DFFSR _14351_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[15]),
    .Q(ALUOut[15]),
    .R(rst_bF$buf29),
    .S(vdd)
);

FILL FILL423320x251940 (
);

FILL FILL88160x345800 (
);

FILL FILL102600x153140 (
);

FILL FILL69920x4940 (
);

FILL FILL_1__16278_ (
);

OR2X2 _15976_ (
    .A(_4922_),
    .B(_4915_),
    .Y(_4923_)
);

OR2X2 _15556_ (
    .A(_4508_),
    .B(_4507_),
    .Y(_4509_)
);

FILL FILL68400x44460 (
);

NOR2X1 _15136_ (
    .A(_4044_),
    .B(_4042_),
    .Y(\datapath_1.regfile_1.regEn [19])
);

AND2X2 _10691_ (
    .A(_1152_),
    .B(_1151_),
    .Y(_1125_[13])
);

AND2X2 _10271_ (
    .A(_932_),
    .B(_931_),
    .Y(_927_[2])
);

FILL FILL_1__8408_ (
);

FILL FILL399000x207480 (
);

FILL FILL_0__16212_ (
);

FILL FILL431680x365560 (
);

FILL FILL266000x296400 (
);

FILL FILL89680x83980 (
);

FILL FILL128440x24700 (
);

FILL FILL_1__12198_ (
);

OR2X2 _11896_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .B(_1784__bF$buf0),
    .Y(_1776_)
);

OR2X2 _11476_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .B(_1586__bF$buf4),
    .Y(_1556_)
);

OR2X2 _11056_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .B(_1388__bF$buf3),
    .Y(_1336_)
);

FILL FILL_0__17837_ (
);

FILL FILL_0__17417_ (
);

AND2X2 _17702_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [5]),
    .Y(_6623_)
);

FILL FILL_0__12972_ (
);

FILL FILL_0__12552_ (
);

FILL FILL_0__12132_ (
);

OR2X2 _9624_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_601_)
);

DFFSR _9204_ (
    .CLK(clk_bF$buf70),
    .D(_333_[6]),
    .Q(\datapath_1.regfile_1.regOut[6] [6]),
    .R(rst_bF$buf66),
    .S(vdd)
);

FILL FILL273600x232180 (
);

AND2X2 _18907_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_7809_)
);

FILL FILL_0__13337_ (
);

AND2X2 _13622_ (
    .A(_3087__bF$buf0),
    .B(\datapath_1.ALUResult [4]),
    .Y(_3113_)
);

AND2X2 _13202_ (
    .A(_2750_),
    .B(_2741_),
    .Y(_2751_)
);

AND2X2 _16094_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_5039_)
);

FILL FILL_0__17590_ (
);

FILL FILL_0__17170_ (
);

FILL FILL_1__15969_ (
);

AND2X2 _14827_ (
    .A(_3917_),
    .B(_3916_),
    .Y(_3870_[23])
);

FILL FILL7600x158080 (
);

AND2X2 _14407_ (
    .A(_3697_),
    .B(_3696_),
    .Y(_3672_[12])
);

INVX1 _17299_ (
    .A(\datapath_1.PCJump [23]),
    .Y(_6225_)
);

FILL FILL_0__15903_ (
);

FILL FILL163400x271700 (
);

FILL FILL463600x54340 (
);

FILL FILL_0__18795_ (
);

OR2X2 _18660_ (
    .A(_7565_),
    .B(_7558_),
    .Y(_7566_)
);

AND2X2 _18240_ (
    .A(_6229__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_7153_)
);

FILL FILL_0__13090_ (
);

FILL FILL_1__11049_ (
);

FILL FILL_0__8896_ (
);

FILL FILL108680x19760 (
);

FILL FILL_0__8476_ (
);

DFFSR _10747_ (
    .CLK(clk_bF$buf34),
    .D(_1125_[1]),
    .Q(\datapath_1.regfile_1.regOut[18] [1]),
    .R(rst_bF$buf71),
    .S(vdd)
);

OR2X2 _10327_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .B(_992__bF$buf2),
    .Y(_970_)
);

FILL FILL_1__12410_ (
);

FILL FILL_0__11823_ (
);

OR2X2 _19445_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_8332_)
);

AND2X2 _19025_ (
    .A(_6323__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_7926_)
);

FILL FILL_0__14295_ (
);

OR2X2 _14580_ (
    .A(memoryOutData[27]),
    .B(_3803__bF$buf1),
    .Y(_3793_)
);

FILL FILL294120x256880 (
);

AND2X2 _14160_ (
    .A(_3551_),
    .B(_3550_),
    .Y(\datapath_1.mux_wd3.dout [5])
);

FILL FILL381520x261820 (
);

FILL FILL91960x311220 (
);

FILL FILL81320x271700 (
);

FILL FILL_1_BUFX2_insert235 (
);

FILL FILL_1_BUFX2_insert237 (
);

FILL FILL_1_BUFX2_insert239 (
);

FILL FILL24320x98800 (
);

FILL FILL319960x19760 (
);

AND2X2 _15785_ (
    .A(_4230__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_4735_)
);

AND2X2 _15365_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_4321_)
);

OR2X2 _10080_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_845_)
);

FILL FILL_0__16861_ (
);

FILL FILL_0__16441_ (
);

FILL FILL394440x39520 (
);

FILL FILL450680x345800 (
);

FILL FILL60800x88920 (
);

DFFSR _11285_ (
    .CLK(clk_bF$buf24),
    .D(_1389_[23]),
    .Q(\datapath_1.regfile_1.regOut[22] [23]),
    .R(rst_bF$buf82),
    .S(vdd)
);

AND2X2 _17931_ (
    .A(_6206__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_6848_)
);

FILL FILL_0__17226_ (
);

AND2X2 _17511_ (
    .A(_6315__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_6435_)
);

FILL FILL57000x306280 (
);

FILL FILL_0__12361_ (
);

FILL FILL207480x0 (
);

FILL FILL291080x54340 (
);

DFFSR _9853_ (
    .CLK(clk_bF$buf107),
    .D(_663_[10]),
    .Q(\datapath_1.regfile_1.regOut[11] [10]),
    .R(rst_bF$buf95),
    .S(vdd)
);

OR2X2 _9433_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .B(_530__bF$buf1),
    .Y(_514_)
);

OR2X2 _9013_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .B(_332__bF$buf1),
    .Y(_294_)
);

FILL FILL28120x98800 (
);

FILL FILL_1__19438_ (
);

AND2X2 _18716_ (
    .A(_6328__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_7621_)
);

FILL FILL_0__13986_ (
);

AND2X2 _13851_ (
    .A(_3300_),
    .B(_3299_),
    .Y(\datapath_1.alu_1.ALUInA [11])
);

FILL FILL_0__13566_ (
);

FILL FILL_0__13146_ (
);

AND2X2 _13431_ (
    .A(_2503_),
    .B(_2156_),
    .Y(_2965_)
);

AND2X2 _13011_ (
    .A(_2570_),
    .B(_2563_),
    .Y(_2571_)
);

FILL FILL255360x0 (
);

OR2X2 _14636_ (
    .A(vdd),
    .B(\datapath_1.a [3]),
    .Y(_3810_)
);

OR2X2 _14216_ (
    .A(\datapath_1.Data [24]),
    .B(_3605__bF$buf4),
    .Y(_3589_)
);

FILL FILL_0__15712_ (
);

FILL FILL_1__19191_ (
);

FILL FILL216600x19760 (
);

FILL FILL_0__18184_ (
);

AND2X2 _10976_ (
    .A(_1302_),
    .B(_1301_),
    .Y(_1257_[22])
);

AND2X2 _10556_ (
    .A(_1082_),
    .B(_1081_),
    .Y(_1059_[11])
);

FILL FILL_1__17504_ (
);

AND2X2 _10136_ (
    .A(_862_),
    .B(_925_),
    .Y(_861_[0])
);

FILL FILL_0__11632_ (
);

FILL FILL_0__11212_ (
);

FILL FILL_0__19389_ (
);

OR2X2 _19254_ (
    .A(_8148_),
    .B(_8150_),
    .Y(_8151_)
);

DFFSR _8704_ (
    .CLK(clk_bF$buf25),
    .D(_69_[22]),
    .Q(\datapath_1.regfile_1.regOut[2] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

FILL FILL_1__13844_ (
);

AND2X2 _12702_ (
    .A(_2265_),
    .B(_2266_),
    .Y(_2267_)
);

FILL FILL_0__12417_ (
);

AND2X2 _15594_ (
    .A(_4154__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_4547_)
);

INVX1 _15174_ (
    .A(\datapath_1.PCJump [18]),
    .Y(_4132_)
);

OR2X2 _9909_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_751_)
);

FILL FILL_0__16670_ (
);

OR2X2 _13907_ (
    .A(\datapath_1.a [30]),
    .B(_3342__bF$buf0),
    .Y(_3338_)
);

FILL FILL324520x34580 (
);

FILL FILL142880x286520 (
);

OR2X2 _16799_ (
    .A(_5731_),
    .B(_5732_),
    .Y(_5733_)
);

AND2X2 _16379_ (
    .A(_4236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_5319_)
);

FILL FILL4560x9880 (
);

OR2X2 _11094_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_1361_)
);

FILL FILL_0__17875_ (
);

FILL FILL483360x281580 (
);

FILL FILL_0__17455_ (
);

AND2X2 _17740_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_6660_)
);

FILL FILL_0__17035_ (
);

AND2X2 _17320_ (
    .A(_6227_),
    .B(_6214_),
    .Y(_6246_)
);

FILL FILL251560x19760 (
);

FILL FILL_0__12590_ (
);

FILL FILL223440x153140 (
);

AND2X2 _9662_ (
    .A(_626_),
    .B(_625_),
    .Y(_597_[14])
);

AND2X2 _9242_ (
    .A(_406_),
    .B(_405_),
    .Y(_399_[3])
);

DFFSR _12299_ (
    .CLK(clk_bF$buf29),
    .D(_1917_[5]),
    .Q(\datapath_1.regfile_1.regOut[30] [5]),
    .R(rst_bF$buf40),
    .S(vdd)
);

OR2X2 _18945_ (
    .A(_7845_),
    .B(_7846_),
    .Y(_7847_)
);

OR2X2 _18525_ (
    .A(_7431_),
    .B(_7432_),
    .Y(_7433_)
);

OR2X2 _18105_ (
    .A(_7016_),
    .B(_7019_),
    .Y(_7020_)
);

FILL FILL_0__13795_ (
);

FILL FILL_0__13375_ (
);

OR2X2 _13660_ (
    .A(_3145_),
    .B(_3142_),
    .Y(\datapath_1.mux_pcsrc.dout [9])
);

XOR2X1 _13240_ (
    .A(_2420_),
    .B(_2744_),
    .Y(_2786_)
);

FILL FILL278920x19760 (
);

FILL FILL462840x19760 (
);

FILL FILL_0__9702_ (
);

FILL FILL212800x296400 (
);

DFFSR _14865_ (
    .CLK(clk_bF$buf58),
    .D(_3870_[13]),
    .Q(_2_[13]),
    .R(rst_bF$buf15),
    .S(vdd)
);

OR2X2 _14445_ (
    .A(memoryOutData[25]),
    .B(_3737__bF$buf2),
    .Y(_3723_)
);

OR2X2 _14025_ (
    .A(_3439_),
    .B(_3440_),
    .Y(_3441_)
);

FILL FILL209760x247000 (
);

FILL FILL_0__15941_ (
);

FILL FILL176320x108680 (
);

FILL FILL394440x232180 (
);

FILL FILL_1__11087_ (
);

OR2X2 _10785_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_1195_)
);

FILL FILL_1__17733_ (
);

DFFSR _10365_ (
    .CLK(clk_bF$buf66),
    .D(_927_[6]),
    .Q(\datapath_1.regfile_1.regOut[15] [6]),
    .R(rst_bF$buf8),
    .S(vdd)
);

FILL FILL_0__16726_ (
);

FILL FILL_0__16306_ (
);

FILL FILL111720x54340 (
);

FILL FILL_0__11861_ (
);

FILL FILL_0__11441_ (
);

FILL FILL427880x237120 (
);

FILL FILL_0__19198_ (
);

AND2X2 _19483_ (
    .A(_8357_),
    .B(_8356_),
    .Y(_8320_[18])
);

OR2X2 _19063_ (
    .A(_7959_),
    .B(_7962_),
    .Y(_7963_)
);

AND2X2 _8933_ (
    .A(_260_),
    .B(_259_),
    .Y(_201_[29])
);

AND2X2 _8513_ (
    .A(_40_),
    .B(_39_),
    .Y(_3_[18])
);

FILL FILL119320x14820 (
);

FILL FILL_0__12646_ (
);

INVX1 _12931_ (
    .A(_2495_),
    .Y(\datapath_1.ALUResult [31])
);

FILL FILL106400x237120 (
);

FILL FILL_0__12226_ (
);

AOI22X1 _12511_ (
    .A(_2105_),
    .B(_2101_),
    .C(_2104_),
    .D(_2102_),
    .Y(RegWrite)
);

FILL FILL_1_BUFX2_insert615 (
);

FILL FILL_1_BUFX2_insert617 (
);

FILL FILL_1_BUFX2_insert619 (
);

FILL FILL212040x311220 (
);

DFFSR _9718_ (
    .CLK(clk_bF$buf79),
    .D(_597_[4]),
    .Q(\datapath_1.regfile_1.regOut[10] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL_1__8675_ (
);

FILL FILL_1__14438_ (
);

FILL FILL_1__14018_ (
);

OR2X2 _13716_ (
    .A(_3193_),
    .B(_3190_),
    .Y(\datapath_1.mux_pcsrc.dout [17])
);

AND2X2 _16188_ (
    .A(_4146__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_5131_)
);

FILL FILL_1__18691_ (
);

FILL FILL_0__17684_ (
);

FILL FILL_0__17264_ (
);

FILL FILL_1__10778_ (
);

FILL FILL_1__10358_ (
);

OR2X2 _9891_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_739_)
);

DFFSR _9471_ (
    .CLK(clk_bF$buf18),
    .D(_465_[15]),
    .Q(\datapath_1.regfile_1.regOut[8] [15]),
    .R(rst_bF$buf107),
    .S(vdd)
);

OR2X2 _9051_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_319_)
);

FILL FILL240920x256880 (
);

FILL FILL_1__19476_ (
);

FILL FILL_1__19056_ (
);

FILL FILL_0__10712_ (
);

OR2X2 _18754_ (
    .A(_7657_),
    .B(_7658_),
    .Y(_7659_)
);

FILL FILL364800x321100 (
);

OR2X2 _18334_ (
    .A(_7244_),
    .B(_7243_),
    .Y(_7245_)
);

FILL FILL_0__18049_ (
);

FILL FILL_0__9931_ (
);

FILL FILL_0__9511_ (
);

FILL FILL_1__15396_ (
);

DFFSR _19539_ (
    .CLK(clk_bF$buf5),
    .D(_8320_[16]),
    .Q(\datapath_1.regfile_1.regOut[0] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

OR2X2 _19119_ (
    .A(_8016_),
    .B(_8017_),
    .Y(_8018_)
);

AND2X2 _14674_ (
    .A(_3835_),
    .B(_3834_),
    .Y(_3804_[15])
);

FILL FILL_0__14389_ (
);

AND2X2 _14254_ (
    .A(_3615_),
    .B(_3614_),
    .Y(_3606_[4])
);

FILL FILL471960x192660 (
);

FILL FILL_0__15330_ (
);

FILL FILL58520x256880 (
);

FILL FILL_1__13709_ (
);

OR2X2 _15879_ (
    .A(_4826_),
    .B(_4825_),
    .Y(_4827_)
);

OR2X2 _15459_ (
    .A(_4413_),
    .B(_4412_),
    .Y(_4414_)
);

OR2X2 _15039_ (
    .A(_4017_),
    .B(_4027_),
    .Y(_4028_)
);

OR2X2 _10594_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_1124__bF$buf1),
    .Y(_1108_)
);

OR2X2 _10174_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .B(_926__bF$buf1),
    .Y(_888_)
);

FILL FILL7600x9880 (
);

FILL FILL_0__16955_ (
);

FILL FILL_0__16535_ (
);

AND2X2 _16820_ (
    .A(_4241__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_5754_)
);

OR2X2 _16400_ (
    .A(_5336_),
    .B(_5339_),
    .Y(_5340_)
);

FILL FILL479560x83980 (
);

FILL FILL158080x14820 (
);

FILL FILL_0__11250_ (
);

OR2X2 _19292_ (
    .A(_8173_),
    .B(_8188_),
    .Y(_8189_)
);

OR2X2 _8742_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_153_)
);

FILL FILL202160x266760 (
);

DFFSR _11799_ (
    .CLK(clk_bF$buf4),
    .D(_1653_[21]),
    .Q(\datapath_1.regfile_1.regOut[26] [21]),
    .R(rst_bF$buf20),
    .S(vdd)
);

OR2X2 _11379_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_1511_)
);

FILL FILL_1__13462_ (
);

AND2X2 _17605_ (
    .A(_6527_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd1 [3])
);

NAND2X1 _12740_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .B(_2304_),
    .Y(_2305_)
);

DFFSR _12320_ (
    .CLK(clk_bF$buf75),
    .D(_1917_[26]),
    .Q(\datapath_1.regfile_1.regOut[30] [26]),
    .R(rst_bF$buf27),
    .S(vdd)
);

FILL FILL365560x133380 (
);

AND2X2 _9947_ (
    .A(_776_),
    .B(_775_),
    .Y(_729_[23])
);

AND2X2 _9527_ (
    .A(_556_),
    .B(_555_),
    .Y(_531_[12])
);

AND2X2 _9107_ (
    .A(_336_),
    .B(_335_),
    .Y(_333_[1])
);

FILL FILL39520x202540 (
);

FILL FILL136800x286520 (
);

FILL FILL19000x88920 (
);

FILL FILL_0_BUFX2_insert270 (
);

FILL FILL_0_BUFX2_insert272 (
);

FILL FILL_0_BUFX2_insert274 (
);

OR2X2 _13945_ (
    .A(_3372_),
    .B(_3369_),
    .Y(\datapath_1.alu_1.ALUInB [3])
);

OR2X2 _13525_ (
    .A(IorD_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [12]),
    .Y(_3038_)
);

OAI21X1 _13105_ (
    .A(_2273_),
    .B(_2376__bF$buf2),
    .C(_2658_),
    .Y(_2659_)
);

FILL FILL_0_BUFX2_insert276 (
);

FILL FILL33440x355680 (
);

FILL FILL438520x247000 (
);

FILL FILL_0_BUFX2_insert278 (
);

FILL FILL_0_BUFX2_insert279 (
);

FILL FILL4560x153140 (
);

FILL FILL_1__18080_ (
);

FILL FILL50920x365560 (
);

FILL FILL_1__10167_ (
);

FILL FILL424080x177840 (
);

OR2X2 _9280_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .B(_464__bF$buf0),
    .Y(_432_)
);

FILL FILL460560x350740 (
);

FILL FILL_0__15806_ (
);

FILL FILL_0__10941_ (
);

FILL FILL_0__18698_ (
);

OR2X2 _18983_ (
    .A(_7883_),
    .B(_7882_),
    .Y(_7884_)
);

AND2X2 _18563_ (
    .A(_6297__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_7471_)
);

FILL FILL_0__18278_ (
);

AND2X2 _18143_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_7057_)
);

FILL FILL_0__8799_ (
);

FILL FILL89680x0 (
);

FILL FILL_0__9320_ (
);

FILL FILL_0__11306_ (
);

OR2X2 _19348_ (
    .A(_8240_),
    .B(_8243_),
    .Y(_8244_)
);

FILL FILL14440x301340 (
);

DFFSR _14483_ (
    .CLK(clk_bF$buf78),
    .D(_3672_[18]),
    .Q(\datapath_1.Data [18]),
    .R(rst_bF$buf110),
    .S(vdd)
);

OR2X2 _14063_ (
    .A(_3473_),
    .B(_3472_),
    .Y(_3474_)
);

FILL FILL318440x212420 (
);

FILL FILL504640x227240 (
);

FILL FILL329840x281580 (
);

FILL FILL344280x153140 (
);

OR2X2 _15688_ (
    .A(_4635_),
    .B(_4638_),
    .Y(_4639_)
);

AND2X2 _15268_ (
    .A(_4225__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_4226_)
);

FILL FILL29640x291460 (
);

FILL FILL_0__16344_ (
);

FILL FILL_1__9901_ (
);

FILL FILL134520x335920 (
);

FILL FILL316160x286520 (
);

DFFSR _8971_ (
    .CLK(clk_bF$buf44),
    .D(_201_[31]),
    .Q(\datapath_1.regfile_1.regOut[4] [31]),
    .R(rst_bF$buf97),
    .S(vdd)
);

OR2X2 _8551_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .B(_68__bF$buf0),
    .Y(_66_)
);

FILL FILL205960x44460 (
);

FILL FILL_1__18556_ (
);

OR2X2 _11188_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .B(_1454__bF$buf1),
    .Y(_1404_)
);

FILL FILL466640x207480 (
);

FILL FILL_0__17549_ (
);

OR2X2 _17834_ (
    .A(_6752_),
    .B(_6751_),
    .Y(_6753_)
);

AND2X2 _17414_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_6339_)
);

FILL FILL_0__17129_ (
);

FILL FILL_0__12684_ (
);

FILL FILL_0__12264_ (
);

OR2X2 _9756_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_669_)
);

DFFSR _9336_ (
    .CLK(clk_bF$buf113),
    .D(_399_[9]),
    .Q(\datapath_1.regfile_1.regOut[7] [9]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL202160x59280 (
);

FILL FILL_1__14896_ (
);

AND2X2 _18619_ (
    .A(_6302__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_7526_)
);

FILL FILL_0__13889_ (
);

FILL FILL_0__13469_ (
);

OR2X2 _13754_ (
    .A(_3224_),
    .B(_3225_),
    .Y(_3226_)
);

AND2X2 _13334_ (
    .A(_2874_),
    .B(_2871_),
    .Y(_2875_)
);

FILL FILL_0__14410_ (
);

FILL FILL223440x316160 (
);

FILL FILL487160x365560 (
);

AND2X2 _14959_ (
    .A(_3985_),
    .B(_3984_),
    .Y(_3936_[24])
);

AND2X2 _14539_ (
    .A(_3765_),
    .B(_3764_),
    .Y(_3738_[13])
);

OR2X2 _14119_ (
    .A(_3521_),
    .B(_3520_),
    .Y(_3522_)
);

FILL FILL_1__16202_ (
);

OR2X2 _15900_ (
    .A(_4846_),
    .B(_4847_),
    .Y(_4848_)
);

FILL FILL_0__10330_ (
);

FILL FILL82080x197600 (
);

AND2X2 _18792_ (
    .A(_6221__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_7696_)
);

OR2X2 _18372_ (
    .A(_7282_),
    .B(_7281_),
    .Y(_7283_)
);

FILL FILL126160x256880 (
);

FILL FILL244720x247000 (
);

DFFSR _10879_ (
    .CLK(clk_bF$buf45),
    .D(_1191_[4]),
    .Q(\datapath_1.regfile_1.regOut[19] [4]),
    .R(rst_bF$buf54),
    .S(vdd)
);

OR2X2 _10459_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_1058__bF$buf1),
    .Y(_1038_)
);

FILL FILL350360x321100 (
);

OR2X2 _10039_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .B(_860__bF$buf1),
    .Y(_818_)
);

FILL FILL_1__12962_ (
);

FILL FILL_1__12542_ (
);

FILL FILL_0__11955_ (
);

OR2X2 _11820_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_1725_)
);

DFFSR _11400_ (
    .CLK(clk_bF$buf102),
    .D(_1455_[9]),
    .Q(\datapath_1.regfile_1.regOut[23] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

AND2X2 _19157_ (
    .A(_6323__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_8056_)
);

OR2X2 _14292_ (
    .A(\datapath_1.ALUResult [17]),
    .B(_3671__bF$buf0),
    .Y(_3641_)
);

OR2X2 _8607_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_83_)
);

INVX1 _12605_ (
    .A(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2170_)
);

OR2X2 _15497_ (
    .A(_4443_),
    .B(_4450_),
    .Y(_4451_)
);

AND2X2 _15077_ (
    .A(_4063_),
    .B(_4041_),
    .Y(_4064_)
);

FILL FILL_0__16993_ (
);

FILL FILL_0__16153_ (
);

FILL FILL107160x202540 (
);

AND2X2 _8780_ (
    .A(_178_),
    .B(_177_),
    .Y(_135_[21])
);

FILL FILL_0__17778_ (
);

OR2X2 _17643_ (
    .A(_6561_),
    .B(_6564_),
    .Y(_6565_)
);

OR2X2 _17223_ (
    .A(_6148_),
    .B(_6149_),
    .Y(_6150_)
);

FILL FILL105640x370500 (
);

FILL FILL127680x83980 (
);

FILL FILL_0__12493_ (
);

FILL FILL_0__12073_ (
);

FILL FILL219640x118560 (
);

DFFSR _9985_ (
    .CLK(clk_bF$buf72),
    .D(_729_[13]),
    .Q(\datapath_1.regfile_1.regOut[12] [13]),
    .R(rst_bF$buf32),
    .S(vdd)
);

OR2X2 _9565_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_596__bF$buf0),
    .Y(_582_)
);

OR2X2 _9145_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .B(_398__bF$buf2),
    .Y(_362_)
);

FILL FILL_0__8400_ (
);

FILL FILL_1__14285_ (
);

AND2X2 _18848_ (
    .A(_6289__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_7751_)
);

FILL FILL_0_BUFX2_insert650 (
);

FILL FILL281960x232180 (
);

NOR2X1 _18428_ (
    .A(_6310__bF$buf2),
    .B(_7337_),
    .Y(_7338_)
);

OR2X2 _18008_ (
    .A(_6923_),
    .B(_6922_),
    .Y(_6924_)
);

FILL FILL_0_BUFX2_insert652 (
);

OR2X2 _13983_ (
    .A(_3403_),
    .B(_3404_),
    .Y(_3405_)
);

FILL FILL_0_BUFX2_insert654 (
);

AND2X2 _13563_ (
    .A(_3063_),
    .B(_3062_),
    .Y(_1_[24])
);

AND2X2 _13143_ (
    .A(_2694_),
    .B(_2686_),
    .Y(_2695_)
);

FILL FILL_0_BUFX2_insert656 (
);

FILL FILL_0_BUFX2_insert658 (
);

FILL FILL_0_BUFX2_insert659 (
);

FILL FILL_0__19504_ (
);

FILL FILL475760x59280 (
);

FILL FILL312360x54340 (
);

FILL FILL409640x375440 (
);

FILL FILL173280x103740 (
);

OR2X2 _14768_ (
    .A(vdd),
    .B(_2_[4]),
    .Y(_3878_)
);

DFFSR _14348_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[12]),
    .Q(ALUOut[12]),
    .R(rst_bF$buf29),
    .S(vdd)
);

FILL FILL_1__16851_ (
);

FILL FILL_0__15844_ (
);

FILL FILL_0__15424_ (
);

FILL FILL291080x321100 (
);

OR2X2 _18181_ (
    .A(_7094_),
    .B(_7093_),
    .Y(_7095_)
);

FILL FILL11400x158080 (
);

FILL FILL334400x232180 (
);

AND2X2 _10688_ (
    .A(_1150_),
    .B(_1149_),
    .Y(_1125_[12])
);

AND2X2 _10268_ (
    .A(_930_),
    .B(_929_),
    .Y(_927_[1])
);

FILL FILL_1__12351_ (
);

FILL FILL_0__16629_ (
);

AND2X2 _16914_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [26]),
    .Y(_5846_)
);

FILL FILL_0__16209_ (
);

FILL FILL_0__11764_ (
);

FILL FILL421040x143260 (
);

FILL FILL231800x83980 (
);

AND2X2 _19386_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_8281_)
);

FILL FILL316160x54340 (
);

FILL FILL338200x153140 (
);

DFFSR _8836_ (
    .CLK(clk_bF$buf81),
    .D(_135_[25]),
    .Q(\datapath_1.regfile_1.regOut[3] [25]),
    .R(rst_bF$buf13),
    .S(vdd)
);

BUFX2 _8416_ (
    .A(_1_[24]),
    .Y(memoryAddress[24])
);

FILL FILL217360x301340 (
);

FILL FILL182400x143260 (
);

FILL FILL_1__13136_ (
);

FILL FILL403560x316160 (
);

FILL FILL_0__12969_ (
);

AND2X2 _12834_ (
    .A(_2398_),
    .B(_2396_),
    .Y(_2399_)
);

FILL FILL_0__12549_ (
);

FILL FILL_0__12129_ (
);

OR2X2 _12414_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_2041_)
);

FILL FILL_0__13910_ (
);

FILL FILL_0__16382_ (
);

FILL FILL121600x14820 (
);

AND2X2 _13619_ (
    .A(_3081__bF$buf1),
    .B(ALUOut[4]),
    .Y(_3110_)
);

FILL FILL251560x227240 (
);

FILL FILL235600x83980 (
);

FILL FILL_1__15702_ (
);

FILL FILL29640x227240 (
);

FILL FILL120080x335920 (
);

FILL FILL_1__18174_ (
);

OR2X2 _17872_ (
    .A(_6786_),
    .B(_6789_),
    .Y(_6790_)
);

AND2X2 _17452_ (
    .A(_6244__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_6377_)
);

FILL FILL_0__17167_ (
);

OR2X2 _17032_ (
    .A(_5961_),
    .B(_5958_),
    .Y(_5962_)
);

AND2X2 _9794_ (
    .A(_694_),
    .B(_693_),
    .Y(_663_[15])
);

AND2X2 _9374_ (
    .A(_474_),
    .B(_473_),
    .Y(_465_[4])
);

FILL FILL_1__11622_ (
);

FILL FILL369360x217360 (
);

DFFSR _10900_ (
    .CLK(clk_bF$buf41),
    .D(_1191_[25]),
    .Q(\datapath_1.regfile_1.regOut[19] [25]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL19760x172900 (
);

FILL FILL490960x29640 (
);

AND2X2 _18657_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_7563_)
);

INVX1 _18237_ (
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_7150_)
);

FILL FILL32680x167960 (
);

OR2X2 _13792_ (
    .A(_3258_),
    .B(_3257_),
    .Y(_3259_)
);

FILL FILL_0__13087_ (
);

NAND3X1 _13372_ (
    .A(_2379__bF$buf3),
    .B(\datapath_1.alu_1.ALUInB [4]),
    .C(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2910_)
);

FILL FILL386840x227240 (
);

FILL FILL_0__19313_ (
);

FILL FILL_1__12827_ (
);

FILL FILL120080x24700 (
);

CLKBUF1 CLKBUF1_insert200 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert201 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert202 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert203 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf20)
);

FILL FILL_0__9834_ (
);

FILL FILL_0__9414_ (
);

CLKBUF1 CLKBUF1_insert204 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert205 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert206 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert207 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert208 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert209 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf14)
);

DFFSR _14997_ (
    .CLK(clk_bF$buf62),
    .D(_3936_[16]),
    .Q(\datapath_1.mux_iord.din0 [16]),
    .R(rst_bF$buf18),
    .S(vdd)
);

OR2X2 _14577_ (
    .A(memoryOutData[26]),
    .B(_3803__bF$buf1),
    .Y(_3791_)
);

AND2X2 _14157_ (
    .A(_3549_),
    .B(_3548_),
    .Y(\datapath_1.mux_wd3.dout [4])
);

FILL FILL_0__15653_ (
);

FILL FILL266000x207480 (
);

FILL FILL402800x167960 (
);

DFFSR _10497_ (
    .CLK(clk_bF$buf51),
    .D(_993_[9]),
    .Q(\datapath_1.regfile_1.regOut[16] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

FILL FILL_1__17025_ (
);

OR2X2 _10077_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_843_)
);

FILL FILL_1__12580_ (
);

FILL FILL_0__16858_ (
);

OR2X2 _16723_ (
    .A(_5656_),
    .B(_5657_),
    .Y(_5658_)
);

FILL FILL_0__16018_ (
);

OR2X2 _16303_ (
    .A(_5241_),
    .B(_5244_),
    .Y(_5245_)
);

FILL FILL_0__11993_ (
);

FILL FILL47120x281580 (
);

FILL FILL_0__11573_ (
);

FILL FILL425600x251940 (
);

AND2X2 _19195_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_8093_)
);

FILL FILL224960x266760 (
);

AND2X2 _8645_ (
    .A(_108_),
    .B(_107_),
    .Y(_69_[19])
);

FILL FILL183920x14820 (
);

FILL FILL_1__13785_ (
);

OR2X2 _17928_ (
    .A(_6814_),
    .B(_6845_),
    .Y(_6846_)
);

AND2X2 _17508_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_6432_)
);

FILL FILL247760x350740 (
);

FILL FILL_0__12778_ (
);

AND2X2 _12643_ (
    .A(_2205_),
    .B(_2207_),
    .Y(_2208_)
);

FILL FILL_0__12358_ (
);

OR2X2 _12223_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .B(_1982__bF$buf2),
    .Y(_1934_)
);

FILL FILL433960x365560 (
);

FILL FILL_0_BUFX2_insert1001 (
);

FILL FILL_0_BUFX2_insert1002 (
);

FILL FILL_0_BUFX2_insert1003 (
);

FILL FILL_0_BUFX2_insert1004 (
);

FILL FILL_0_BUFX2_insert1005 (
);

FILL FILL_0_BUFX2_insert1007 (
);

FILL FILL3800x167960 (
);

FILL FILL_0_BUFX2_insert1009 (
);

AND2X2 _13848_ (
    .A(_3298_),
    .B(_3297_),
    .Y(\datapath_1.alu_1.ALUInA [10])
);

AND2X2 _13428_ (
    .A(_2956_),
    .B(_2962_),
    .Y(_2963_)
);

XOR2X1 _13008_ (
    .A(_2540_),
    .B(_2556_),
    .Y(_2568_)
);

FILL FILL_0__14504_ (
);

FILL FILL_0__17396_ (
);

INVX1 _17681_ (
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_6602_)
);

AND2X2 _17261_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_6188_)
);

FILL FILL345040x133380 (
);

FILL FILL_1__16716_ (
);

OR2X2 _9183_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_387_)
);

FILL FILL_0__15709_ (
);

FILL FILL_0__10844_ (
);

FILL FILL49400x74100 (
);

FILL FILL_0__10004_ (
);

AND2X2 _18886_ (
    .A(_6287__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_7789_)
);

AND2X2 _18466_ (
    .A(_6247__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_7375_)
);

AND2X2 _18046_ (
    .A(_6238__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_6962_)
);

AND2X2 _13181_ (
    .A(_2729_),
    .B(_2242_),
    .Y(_2730_)
);

FILL FILL161880x158080 (
);

FILL FILL342000x93860 (
);

FILL FILL148200x261820 (
);

FILL FILL_0__9643_ (
);

DFFSR _11914_ (
    .CLK(clk_bF$buf54),
    .D(_1719_[7]),
    .Q(\datapath_1.regfile_1.regOut[27] [7]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL_0__11209_ (
);

FILL FILL245480x212420 (
);

AND2X2 _14386_ (
    .A(_3683_),
    .B(_3682_),
    .Y(_3672_[5])
);

FILL FILL_0__15882_ (
);

FILL FILL_0__15462_ (
);

FILL FILL_0__15042_ (
);

FILL FILL363280x0 (
);

FILL FILL171000x83980 (
);

FILL FILL_1__17674_ (
);

OR2X2 _16952_ (
    .A(_5883_),
    .B(_5868_),
    .Y(_5884_)
);

AND2X2 _16532_ (
    .A(_4181__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_5470_)
);

FILL FILL_0__16247_ (
);

AND2X2 _16112_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_5057_)
);

FILL FILL296400x256880 (
);

FILL FILL_0__11382_ (
);

FILL FILL370880x98800 (
);

OR2X2 _8874_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_221_)
);

BUFX2 _8454_ (
    .A(_2_[30]),
    .Y(memoryWriteData[30])
);

FILL FILL_1__18039_ (
);

AND2X2 _17737_ (
    .A(_6232__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_6657_)
);

AND2X2 _17317_ (
    .A(_6219_),
    .B(_6214_),
    .Y(_6243_)
);

NAND3X1 _12872_ (
    .A(_2436_),
    .B(\datapath_1.alu_1.ALUInB [10]),
    .C(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2437_)
);

DFFSR _12452_ (
    .CLK(clk_bF$buf78),
    .D(_1983_[29]),
    .Q(\datapath_1.regfile_1.regOut[31] [29]),
    .R(rst_bF$buf110),
    .S(vdd)
);

AND2X2 _12032_ (
    .A(_1846_),
    .B(_1845_),
    .Y(_1785_[30])
);

FILL FILL_0__18813_ (
);

AND2X2 _9659_ (
    .A(_624_),
    .B(_623_),
    .Y(_597_[13])
);

AND2X2 _9239_ (
    .A(_404_),
    .B(_403_),
    .Y(_399_[2])
);

FILL FILL_0__8914_ (
);

AND2X2 _13657_ (
    .A(_3087__bF$buf1),
    .B(\datapath_1.ALUResult [9]),
    .Y(_3143_)
);

NOR2X1 _13237_ (
    .A(_2503_),
    .B(_2215_),
    .Y(_2783_)
);

FILL FILL_1__15320_ (
);

OR2X2 _17490_ (
    .A(_6413_),
    .B(_6409_),
    .Y(_6414_)
);

OR2X2 _17070_ (
    .A(_5999_),
    .B(_5998_),
    .Y(_6000_)
);

FILL FILL273600x74100 (
);

FILL FILL290320x24700 (
);

FILL FILL_1__16525_ (
);

FILL FILL389120x158080 (
);

FILL FILL_1__11240_ (
);

FILL FILL_0__15518_ (
);

AND2X2 _15803_ (
    .A(_4241__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_4752_)
);

FILL FILL_0__10653_ (
);

FILL FILL505400x345800 (
);

AND2X2 _18695_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_7601_)
);

OR2X2 _18275_ (
    .A(_7183_),
    .B(_7186_),
    .Y(_7187_)
);

FILL FILL275120x276640 (
);

AND2X2 _11723_ (
    .A(_1680_),
    .B(_1679_),
    .Y(_1653_[13])
);

FILL FILL_0__9032_ (
);

AND2X2 _11303_ (
    .A(_1460_),
    .B(_1459_),
    .Y(_1455_[2])
);

FILL FILL22800x29640 (
);

OR2X2 _14195_ (
    .A(\datapath_1.Data [17]),
    .B(_3605__bF$buf2),
    .Y(_3575_)
);

FILL FILL423320x19760 (
);

FILL FILL129960x39520 (
);

FILL FILL_0__15271_ (
);

FILL FILL66880x256880 (
);

FILL FILL_1_BUFX2_insert580 (
);

OR2X2 _12928_ (
    .A(_2387__bF$buf2),
    .B(_2492_),
    .Y(_2493_)
);

FILL FILL_1_BUFX2_insert582 (
);

FILL FILL493240x266760 (
);

NAND3X1 _12508_ (
    .A(_2103_),
    .B(\control_1.reg_state.dout [2]),
    .C(_2100_),
    .Y(_2104_)
);

FILL FILL_1__17063_ (
);

FILL FILL_0__16896_ (
);

OR2X2 _16761_ (
    .A(_5695_),
    .B(_5664_),
    .Y(_5696_)
);

FILL FILL_0__16476_ (
);

AND2X2 _16341_ (
    .A(_4210__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_5282_)
);

FILL FILL_0__11191_ (
);

DFFSR _8683_ (
    .CLK(clk_bF$buf43),
    .D(_69_[1]),
    .Q(\datapath_1.regfile_1.regOut[2] [1]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL256120x222300 (
);

FILL FILL_1__10931_ (
);

BUFX2 BUFX2_insert250 (
    .A(_4146_),
    .Y(_4146__bF$buf3)
);

BUFX2 BUFX2_insert251 (
    .A(_4146_),
    .Y(_4146__bF$buf2)
);

BUFX2 BUFX2_insert252 (
    .A(_4146_),
    .Y(_4146__bF$buf1)
);

BUFX2 BUFX2_insert253 (
    .A(_4146_),
    .Y(_4146__bF$buf0)
);

OR2X2 _17966_ (
    .A(_6881_),
    .B(_6882_),
    .Y(_6883_)
);

BUFX2 BUFX2_insert254 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf4 )
);

OR2X2 _17546_ (
    .A(_6467_),
    .B(_6468_),
    .Y(_6469_)
);

BUFX2 BUFX2_insert255 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf3 )
);

BUFX2 BUFX2_insert256 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf2 )
);

OR2X2 _17126_ (
    .A(_6054_),
    .B(_6053_),
    .Y(_6055_)
);

BUFX2 BUFX2_insert257 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf1 )
);

BUFX2 BUFX2_insert258 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf0 )
);

FILL FILL_0__12396_ (
);

BUFX2 BUFX2_insert259 (
    .A(_6271_),
    .Y(_6271__bF$buf4)
);

XOR2X1 _12681_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2246_)
);

OR2X2 _12261_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[30] [21]),
    .Y(_1959_)
);

FILL FILL_0__18622_ (
);

FILL FILL127680x276640 (
);

OR2X2 _9888_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_737_)
);

DFFSR _9468_ (
    .CLK(clk_bF$buf102),
    .D(_465_[12]),
    .Q(\datapath_1.regfile_1.regOut[8] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

OR2X2 _9048_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_317_)
);

FILL FILL_0__8723_ (
);

OR2X2 _13886_ (
    .A(\datapath_1.a [23]),
    .B(_3342__bF$buf4),
    .Y(_3324_)
);

AND2X2 _13466_ (
    .A(_2986_),
    .B(_2998_),
    .Y(_2999_)
);

AND2X2 _13046_ (
    .A(_2602_),
    .B(_2308_),
    .Y(_2603_)
);

FILL FILL307040x9880 (
);

FILL FILL_0__19407_ (
);

FILL FILL_0__14122_ (
);

FILL FILL212800x207480 (
);

FILL FILL113240x103740 (
);

FILL FILL_0__9928_ (
);

FILL FILL130720x113620 (
);

FILL FILL_0__15747_ (
);

FILL FILL266760x0 (
);

FILL FILL_0__15327_ (
);

AND2X2 _15612_ (
    .A(_4154__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_4564_)
);

FILL FILL_0__10462_ (
);

FILL FILL_0__10042_ (
);

OR2X2 _18084_ (
    .A(_6998_),
    .B(_6997_),
    .Y(_6999_)
);

FILL FILL329840x4940 (
);

FILL FILL365560x9880 (
);

FILL FILL_0__19160_ (
);

FILL FILL_1__17539_ (
);

AND2X2 _16817_ (
    .A(_4236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_5751_)
);

FILL FILL504640x113620 (
);

FILL FILL278160x19760 (
);

OR2X2 _11952_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_1793_)
);

FILL FILL_0__9261_ (
);

DFFSR _11532_ (
    .CLK(clk_bF$buf28),
    .D(_1521_[12]),
    .Q(\datapath_1.regfile_1.regOut[24] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

FILL FILL_0__11247_ (
);

OR2X2 _11112_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_1373_)
);

OR2X2 _19289_ (
    .A(_8185_),
    .B(_8184_),
    .Y(_8186_)
);

FILL FILL348840x4940 (
);

OR2X2 _8739_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_151_)
);

FILL FILL178600x108680 (
);

FILL FILL_1__13879_ (
);

FILL FILL328320x4940 (
);

FILL FILL151240x271700 (
);

FILL FILL79040x232180 (
);

FILL FILL198360x34580 (
);

AND2X2 _12737_ (
    .A(_2295_),
    .B(_2301_),
    .Y(_2302_)
);

DFFSR _12317_ (
    .CLK(clk_bF$buf101),
    .D(_1917_[23]),
    .Q(\datapath_1.regfile_1.regOut[30] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL_0__13813_ (
);

FILL FILL_1__17292_ (
);

AND2X2 _16990_ (
    .A(_4135__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_5921_)
);

AND2X2 _16570_ (
    .A(_5507_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [20])
);

FILL FILL_0__16285_ (
);

OR2X2 _16150_ (
    .A(_5092_),
    .B(_5093_),
    .Y(_5094_)
);

AND2X2 _8492_ (
    .A(_26_),
    .B(_25_),
    .Y(_3_[11])
);

FILL FILL_1__10320_ (
);

FILL FILL_1__18497_ (
);

FILL FILL199120x266760 (
);

FILL FILL420280x49400 (
);

AND2X2 _17775_ (
    .A(_6221__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_6695_)
);

AND2X2 _17355_ (
    .A(_6280_),
    .B(_6277_),
    .Y(_6281_)
);

FILL FILL286520x271700 (
);

FILL FILL214320x311220 (
);

NOR2X1 _12490_ (
    .A(_2094_),
    .B(_2091_),
    .Y(BranchNe)
);

OR2X2 _12070_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(_1916__bF$buf4),
    .Y(_1852_)
);

FILL FILL_0__18431_ (
);

FILL FILL_0__18011_ (
);

OR2X2 _9697_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .B(_662__bF$buf4),
    .Y(_650_)
);

OR2X2 _9277_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .B(_464__bF$buf3),
    .Y(_430_)
);

FILL FILL309320x217360 (
);

FILL FILL119320x88920 (
);

FILL FILL_0__8532_ (
);

FILL FILL_0__10938_ (
);

OR2X2 _10803_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_1207_)
);

OR2X2 _13695_ (
    .A(_3175_),
    .B(_3172_),
    .Y(\datapath_1.mux_pcsrc.dout [14])
);

AND2X2 _13275_ (
    .A(_2818_),
    .B(_2809_),
    .Y(_2819_)
);

AND2X2 _19501_ (
    .A(_8369_),
    .B(_8368_),
    .Y(_8320_[24])
);

FILL FILL240160x118560 (
);

FILL FILL_0__9317_ (
);

FILL FILL_1__16143_ (
);

FILL FILL_0__15976_ (
);

AND2X2 _15841_ (
    .A(_4208__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_4790_)
);

FILL FILL_0__15136_ (
);

OR2X2 _15421_ (
    .A(_4374_),
    .B(_4375_),
    .Y(_4376_)
);

DFFSR _15001_ (
    .CLK(clk_bF$buf62),
    .D(_3936_[20]),
    .Q(\datapath_1.mux_iord.din0 [20]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL_0__10691_ (
);

FILL FILL_0__10271_ (
);

FILL FILL344280x64220 (
);

FILL FILL375440x118560 (
);

OR2X2 _16626_ (
    .A(_5561_),
    .B(_5562_),
    .Y(_5563_)
);

AND2X2 _16206_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_5149_)
);

FILL FILL_0__11896_ (
);

OR2X2 _11761_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .B(_1718__bF$buf4),
    .Y(_1706_)
);

OR2X2 _11341_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .B(_1520__bF$buf2),
    .Y(_1486_)
);

FILL FILL_0__11056_ (
);

OR2X2 _19098_ (
    .A(_7966_),
    .B(_7997_),
    .Y(_7998_)
);

FILL FILL_0__17702_ (
);

DFFSR _8968_ (
    .CLK(clk_bF$buf91),
    .D(_201_[28]),
    .Q(\datapath_1.regfile_1.regOut[4] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

OR2X2 _8548_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .B(_68__bF$buf3),
    .Y(_64_)
);

FILL FILL_1__13268_ (
);

FILL FILL_1_BUFX2_insert960 (
);

FILL FILL_1_BUFX2_insert962 (
);

INVX1 _12966_ (
    .A(_2528_),
    .Y(\datapath_1.ALUResult [29])
);

AND2X2 _12546_ (
    .A(_2134_),
    .B(_2120_),
    .Y(_2135_)
);

OR2X2 _12126_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_1889_)
);

FILL FILL_0__18907_ (
);

FILL FILL_0__13622_ (
);

FILL FILL_0__13202_ (
);

FILL FILL_0__16094_ (
);

FILL FILL_1__9651_ (
);

FILL FILL411160x321100 (
);

FILL FILL_0__14827_ (
);

FILL FILL_0__14407_ (
);

BUFX2 BUFX2_insert630 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf9)
);

BUFX2 BUFX2_insert631 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf8)
);

BUFX2 BUFX2_insert632 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf7)
);

BUFX2 BUFX2_insert633 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf6)
);

BUFX2 BUFX2_insert634 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf5)
);

BUFX2 BUFX2_insert635 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf4)
);

OR2X2 _17584_ (
    .A(_6505_),
    .B(_6506_),
    .Y(_6507_)
);

FILL FILL_0__17299_ (
);

BUFX2 BUFX2_insert636 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf3)
);

OR2X2 _17164_ (
    .A(_6091_),
    .B(_6090_),
    .Y(_6092_)
);

FILL FILL227240x350740 (
);

FILL FILL53200x182780 (
);

BUFX2 BUFX2_insert637 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf2)
);

BUFX2 BUFX2_insert638 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf1)
);

BUFX2 BUFX2_insert639 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf0)
);

FILL FILL_0__18660_ (
);

FILL FILL368600x9880 (
);

FILL FILL253080x291460 (
);

FILL FILL_1__16619_ (
);

DFFSR _9086_ (
    .CLK(clk_bF$buf6),
    .D(_267_[17]),
    .Q(\datapath_1.regfile_1.regOut[5] [17]),
    .R(rst_bF$buf6),
    .S(vdd)
);

FILL FILL67640x143260 (
);

FILL FILL_0__8761_ (
);

FILL FILL35720x355680 (
);

FILL FILL_0__10327_ (
);

OR2X2 _10612_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_1124__bF$buf3),
    .Y(_1120_)
);

OR2X2 _18789_ (
    .A(_7689_),
    .B(_7692_),
    .Y(_7693_)
);

OR2X2 _18369_ (
    .A(_7278_),
    .B(_7279_),
    .Y(_7280_)
);

OR2X2 _13084_ (
    .A(_2387__bF$buf1),
    .B(_2638_),
    .Y(_2639_)
);

FILL FILL_0__19445_ (
);

FILL FILL_0__19025_ (
);

OR2X2 _19310_ (
    .A(_8202_),
    .B(_8205_),
    .Y(_8206_)
);

FILL FILL_0__14580_ (
);

FILL FILL426360x177840 (
);

FILL FILL_0__9966_ (
);

FILL FILL_0__9546_ (
);

FILL FILL_0__9126_ (
);

OR2X2 _11817_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_1723_)
);

OR2X2 _14289_ (
    .A(\datapath_1.ALUResult [16]),
    .B(_3671__bF$buf0),
    .Y(_3639_)
);

FILL FILL_1__16792_ (
);

FILL FILL_0__15365_ (
);

AND2X2 _15650_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_4602_)
);

AND2X2 _15230_ (
    .A(_4187__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_4188_)
);

FILL FILL_0__10080_ (
);

FILL FILL_1__8922_ (
);

FILL FILL128440x163020 (
);

FILL FILL_1__17157_ (
);

FILL FILL_1__12292_ (
);

OR2X2 _16855_ (
    .A(_5784_),
    .B(_5787_),
    .Y(_5788_)
);

AND2X2 _16435_ (
    .A(_4230__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_5375_)
);

OR2X2 _16015_ (
    .A(_4959_),
    .B(_4960_),
    .Y(_4961_)
);

AND2X2 _11990_ (
    .A(_1818_),
    .B(_1817_),
    .Y(_1785_[16])
);

AND2X2 _11570_ (
    .A(_1598_),
    .B(_1597_),
    .Y(_1587_[5])
);

DFFSR _11150_ (
    .CLK(clk_bF$buf64),
    .D(_1323_[17]),
    .Q(\datapath_1.regfile_1.regOut[21] [17]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL433960x0 (
);

FILL FILL_0__17931_ (
);

FILL FILL_0__17511_ (
);

FILL FILL42560x242060 (
);

AND2X2 _8777_ (
    .A(_176_),
    .B(_175_),
    .Y(_135_[20])
);

INVX1 _12775_ (
    .A(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2340_)
);

OR2X2 _12355_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .B(_2048__bF$buf2),
    .Y(_2002_)
);

FILL FILL_1__19303_ (
);

FILL FILL_0__13851_ (
);

FILL FILL_0__13011_ (
);

FILL FILL136800x335920 (
);

FILL FILL181640x118560 (
);

FILL FILL_1__9040_ (
);

FILL FILL228760x44460 (
);

FILL FILL_1__15643_ (
);

FILL FILL405080x197600 (
);

FILL FILL266000x88920 (
);

FILL FILL19760x14820 (
);

FILL FILL_0__14636_ (
);

OR2X2 _14921_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [12]),
    .Y(_3960_)
);

OR2X2 _14501_ (
    .A(IRWrite_bF$buf0),
    .B(\aluControl_1.inst [1]),
    .Y(_3740_)
);

FILL FILL_0__14216_ (
);

FILL FILL441560x370500 (
);

OR2X2 _17393_ (
    .A(_6318_),
    .B(_6316_),
    .Y(_6319_)
);

FILL FILL8360x123500 (
);

FILL FILL304000x113620 (
);

FILL FILL_1__16008_ (
);

FILL FILL_1__11983_ (
);

AND2X2 _15706_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [7]),
    .Y(_4657_)
);

FILL FILL86640x123500 (
);

FILL FILL_0__10976_ (
);

AND2X2 _10841_ (
    .A(_1232_),
    .B(_1231_),
    .Y(_1191_[20])
);

AND2X2 _10421_ (
    .A(_1012_),
    .B(_1011_),
    .Y(_993_[9])
);

FILL FILL_0__10136_ (
);

DFFSR _10001_ (
    .CLK(clk_bF$buf88),
    .D(_729_[29]),
    .Q(\datapath_1.regfile_1.regOut[12] [29]),
    .R(rst_bF$buf95),
    .S(vdd)
);

NOR2X1 _18598_ (
    .A(_6310__bF$buf2),
    .B(_7504_),
    .Y(_7505_)
);

INVX1 _18178_ (
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_7092_)
);

FILL FILL367080x177840 (
);

FILL FILL_0__19254_ (
);

FILL FILL_1__12768_ (
);

FILL FILL_0__9775_ (
);

OR2X2 _11626_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .B(_1652__bF$buf4),
    .Y(_1636_)
);

OR2X2 _11206_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .B(_1454__bF$buf2),
    .Y(_1416_)
);

OR2X2 _14098_ (
    .A(_3503_),
    .B(_3502_),
    .Y(_3504_)
);

FILL FILL335160x311220 (
);

FILL FILL_0__15594_ (
);

FILL FILL_1__8731_ (
);

FILL FILL352640x321100 (
);

FILL FILL_0__13907_ (
);

FILL FILL499320x98800 (
);

FILL FILL_0__16799_ (
);

OR2X2 _16664_ (
    .A(_5592_),
    .B(_5599_),
    .Y(_5600_)
);

AND2X2 _16244_ (
    .A(_4135__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_5187_)
);

FILL FILL_0__11094_ (
);

FILL FILL_1__9936_ (
);

FILL FILL_0__17740_ (
);

FILL FILL91960x133380 (
);

INVX2 _8586_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .Y(_134_)
);

FILL FILL458280x69160 (
);

AND2X2 _17869_ (
    .A(_6259__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_6787_)
);

AND2X2 _17449_ (
    .A(_6289__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_6374_)
);

AND2X2 _17029_ (
    .A(_4187__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_5959_)
);

FILL FILL411160x39520 (
);

DFFSR _12584_ (
    .CLK(clk_bF$buf20),
    .D(_2143_[0]),
    .Q(\control_1.reg_state.dout [0]),
    .R(rst_bF$buf22),
    .S(vdd)
);

AND2X2 _12164_ (
    .A(_1914_),
    .B(_1913_),
    .Y(_1851_[31])
);

AND2X2 _18810_ (
    .A(_6255__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_7714_)
);

FILL FILL_0__18525_ (
);

FILL FILL_0__18105_ (
);

FILL FILL_0__13660_ (
);

FILL FILL_0__13240_ (
);

FILL FILL450680x167960 (
);

FILL FILL_0__8626_ (
);

OR2X2 _13789_ (
    .A(_3254_),
    .B(_3255_),
    .Y(_3256_)
);

NAND2X1 _13369_ (
    .A(_2524_),
    .B(_2906_),
    .Y(_2907_)
);

FILL FILL418760x24700 (
);

DFFSR _14730_ (
    .CLK(clk_bF$buf15),
    .D(_3804_[7]),
    .Q(\datapath_1.a [7]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL_0__14445_ (
);

OR2X2 _14310_ (
    .A(\datapath_1.ALUResult [23]),
    .B(_3671__bF$buf1),
    .Y(_3653_)
);

FILL FILL107920x370500 (
);

FILL FILL373160x345800 (
);

FILL FILL120840x365560 (
);

CLKBUF1 CLKBUF1_insert170 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert171 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert172 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert173 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert174 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert175 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert176 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert177 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert178 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert179 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf44)
);

FILL FILL240920x4940 (
);

FILL FILL262200x123500 (
);

FILL FILL_1__16657_ (
);

FILL FILL_1__11372_ (
);

AND2X2 _15935_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_4882_)
);

AND2X2 _15515_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [4]),
    .Y(_4469_)
);

FILL FILL160360x44460 (
);

FILL FILL_0__10785_ (
);

INVX2 _10650_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .Y(_1190_)
);

DFFSR _10230_ (
    .CLK(clk_bF$buf96),
    .D(_861_[0]),
    .Q(\datapath_1.regfile_1.regOut[14] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL_0__19483_ (
);

FILL FILL_0__19063_ (
);

FILL FILL431680x113620 (
);

FILL FILL175560x103740 (
);

FILL FILL_1__12997_ (
);

FILL FILL_1__18803_ (
);

AND2X2 _11855_ (
    .A(_1748_),
    .B(_1747_),
    .Y(_1719_[14])
);

FILL FILL_0__9164_ (
);

AND2X2 _11435_ (
    .A(_1528_),
    .B(_1527_),
    .Y(_1521_[3])
);

DFFSR _11015_ (
    .CLK(clk_bF$buf73),
    .D(_1257_[11]),
    .Q(\datapath_1.regfile_1.regOut[20] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL_0__12931_ (
);

FILL FILL_0__12511_ (
);

FILL FILL342760x276640 (
);

FILL FILL348080x350740 (
);

FILL FILL187720x44460 (
);

FILL FILL371640x44460 (
);

FILL FILL259920x286520 (
);

FILL FILL19000x232180 (
);

FILL FILL_0__13716_ (
);

FILL FILL423320x143260 (
);

FILL FILL167200x133380 (
);

OR2X2 _16893_ (
    .A(_5823_),
    .B(_5824_),
    .Y(_5825_)
);

OR2X2 _16473_ (
    .A(_5396_),
    .B(_5411_),
    .Y(_5412_)
);

FILL FILL_0__16188_ (
);

OR2X2 _16053_ (
    .A(_4997_),
    .B(_4998_),
    .Y(_4999_)
);

FILL FILL_1__9325_ (
);

FILL FILL323000x237120 (
);

FILL FILL231040x83980 (
);

FILL FILL_1__15508_ (
);

BUFX2 _8395_ (
    .A(_1_[3]),
    .Y(memoryAddress[3])
);

FILL FILL446880x9880 (
);

FILL FILL405840x316160 (
);

AND2X2 _17678_ (
    .A(_6229__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_6599_)
);

AND2X2 _17258_ (
    .A(_4130__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_6185_)
);

OR2X2 _12393_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_2027_)
);

FILL FILL190000x311220 (
);

FILL FILL317680x281580 (
);

FILL FILL_0__18754_ (
);

FILL FILL236360x217360 (
);

FILL FILL_1__11428_ (
);

FILL FILL_0__8855_ (
);

AND2X2 _10706_ (
    .A(_1162_),
    .B(_1161_),
    .Y(_1125_[18])
);

FILL FILL253840x227240 (
);

FILL FILL76760x49400 (
);

FILL FILL319200x24700 (
);

AND2X2 _13598_ (
    .A(_3081__bF$buf0),
    .B(ALUOut[1]),
    .Y(_3092_)
);

INVX1 _13178_ (
    .A(_2727_),
    .Y(\datapath_1.ALUResult [16])
);

FILL FILL_1__15261_ (
);

OR2X2 _19404_ (
    .A(_8298_),
    .B(_8297_),
    .Y(_8299_)
);

FILL FILL_0__19119_ (
);

FILL FILL_0__14254_ (
);

FILL FILL121600x88920 (
);

FILL FILL53960x330980 (
);

FILL FILL_1__11181_ (
);

FILL FILL_0__15879_ (
);

FILL FILL34960x167960 (
);

OR2X2 _15744_ (
    .A(_4692_),
    .B(_4693_),
    .Y(_4694_)
);

FILL FILL_0__15459_ (
);

OR2X2 _15324_ (
    .A(_4279_),
    .B(_4280_),
    .Y(_4281_)
);

FILL FILL_0__10594_ (
);

FILL FILL458280x128440 (
);

FILL FILL_0__16820_ (
);

FILL FILL_0__16400_ (
);

FILL FILL114000x365560 (
);

OR2X2 _16949_ (
    .A(_5880_),
    .B(_5879_),
    .Y(_5881_)
);

AND2X2 _16529_ (
    .A(_4234__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_5467_)
);

AND2X2 _16109_ (
    .A(_4175__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_5054_)
);

FILL FILL_0__9393_ (
);

FILL FILL_0__11379_ (
);

DFFSR _11664_ (
    .CLK(clk_bF$buf39),
    .D(_1587_[15]),
    .Q(\datapath_1.regfile_1.regOut[25] [15]),
    .R(rst_bF$buf3),
    .S(vdd)
);

OR2X2 _11244_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_1441_)
);

FILL FILL_0__17605_ (
);

FILL FILL_0__12740_ (
);

AND2X2 _9812_ (
    .A(_706_),
    .B(_705_),
    .Y(_663_[21])
);

OR2X2 _12869_ (
    .A(_2427_),
    .B(_2433_),
    .Y(_2434_)
);

DFFSR _12449_ (
    .CLK(clk_bF$buf55),
    .D(_1983_[26]),
    .Q(\datapath_1.regfile_1.regOut[31] [26]),
    .R(rst_bF$buf24),
    .S(vdd)
);

FILL FILL182400x79040 (
);

AND2X2 _12029_ (
    .A(_1844_),
    .B(_1843_),
    .Y(_1785_[29])
);

FILL FILL_1__14112_ (
);

OR2X2 _13810_ (
    .A(_3272_),
    .B(_3273_),
    .Y(_3274_)
);

FILL FILL_0__13105_ (
);

AND2X2 _16282_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_5224_)
);

FILL FILL332880x340860 (
);

FILL FILL_1__15737_ (
);

FILL FILL_1__10452_ (
);

NOR2X1 _17487_ (
    .A(_6310__bF$buf0),
    .B(_6410_),
    .Y(_6411_)
);

OR2X2 _17067_ (
    .A(_5996_),
    .B(_5995_),
    .Y(_5997_)
);

FILL FILL275880x291460 (
);

FILL FILL_0__18563_ (
);

FILL FILL_0__18143_ (
);

FILL FILL473480x321100 (
);

FILL FILL_0__8664_ (
);

OR2X2 _10935_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_1275_)
);

DFFSR _10515_ (
    .CLK(clk_bF$buf70),
    .D(_993_[27]),
    .Q(\datapath_1.regfile_1.regOut[16] [27]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL198360x148200 (
);

FILL FILL_0__19348_ (
);

NOR2X1 _19213_ (
    .A(_6310__bF$buf1),
    .B(_8110_),
    .Y(_8111_)
);

FILL FILL_0__14063_ (
);

FILL FILL142880x59280 (
);

FILL FILL_0__9449_ (
);

FILL FILL347320x133380 (
);

FILL FILL60800x232180 (
);

AND2X2 _15973_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_4920_)
);

FILL FILL_0__15688_ (
);

FILL FILL_0__15268_ (
);

OR2X2 _15553_ (
    .A(_4505_),
    .B(_4502_),
    .Y(_4506_)
);

NAND2X1 _15133_ (
    .A(_4024_),
    .B(_4009_),
    .Y(_4106_)
);

OR2X2 _16758_ (
    .A(_5689_),
    .B(_5692_),
    .Y(_5693_)
);

AND2X2 _16338_ (
    .A(_4172__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_5279_)
);

OR2X2 _11893_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .B(_1784__bF$buf1),
    .Y(_1774_)
);

FILL FILL_0__11188_ (
);

FILL FILL_1__18421_ (
);

OR2X2 _11473_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .B(_1586__bF$buf4),
    .Y(_1554_)
);

OR2X2 _11053_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .B(_1388__bF$buf3),
    .Y(_1334_)
);

FILL FILL228760x370500 (
);

OR2X2 _9621_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_599_)
);

DFFSR _9201_ (
    .CLK(clk_bF$buf56),
    .D(_333_[3]),
    .Q(\datapath_1.regfile_1.regOut[6] [3]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL45600x177840 (
);

OR2X2 _12678_ (
    .A(_2217_),
    .B(_2242_),
    .Y(_2243_)
);

OR2X2 _12258_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_1957_)
);

OR2X2 _18904_ (
    .A(_7772_),
    .B(_7806_),
    .Y(_7807_)
);

FILL FILL_0__18619_ (
);

FILL FILL465880x34580 (
);

FILL FILL_0__13754_ (
);

FILL FILL_0__13334_ (
);

FILL FILL202920x182780 (
);

AND2X2 _16091_ (
    .A(_4200__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_5036_)
);

FILL FILL239400x242060 (
);

FILL FILL395960x207480 (
);

FILL FILL_1__9783_ (
);

FILL FILL_1__15126_ (
);

FILL FILL_0__14959_ (
);

AND2X2 _14824_ (
    .A(_3915_),
    .B(_3914_),
    .Y(_3870_[22])
);

FILL FILL_0__14539_ (
);

FILL FILL_0__14119_ (
);

AND2X2 _14404_ (
    .A(_3695_),
    .B(_3694_),
    .Y(_3672_[11])
);

AND2X2 _17296_ (
    .A(_6221__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_6222_)
);

FILL FILL_0__15900_ (
);

FILL FILL_0__18792_ (
);

FILL FILL_0__18372_ (
);

OR2X2 _15609_ (
    .A(_4561_),
    .B(_4530_),
    .Y(_4562_)
);

FILL FILL_0__8893_ (
);

FILL FILL_0__8473_ (
);

OR2X2 _10744_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .B(_1190__bF$buf2),
    .Y(_1188_)
);

FILL FILL_0__10039_ (
);

OR2X2 _10324_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .B(_992__bF$buf0),
    .Y(_968_)
);

FILL FILL_0__11820_ (
);

OR2X2 _19442_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_8330_)
);

OR2X2 _19022_ (
    .A(_7922_),
    .B(_7921_),
    .Y(_7923_)
);

FILL FILL_0__14292_ (
);

FILL FILL_0__9678_ (
);

OR2X2 _11949_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[28] [3]),
    .Y(_1791_)
);

FILL FILL_0__9258_ (
);

DFFSR _11529_ (
    .CLK(clk_bF$buf113),
    .D(_1521_[9]),
    .Q(\datapath_1.regfile_1.regOut[24] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

OR2X2 _11109_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_1371_)
);

FILL FILL_0__12605_ (
);

FILL FILL_1__16084_ (
);

OR2X2 _15782_ (
    .A(_4730_),
    .B(_4731_),
    .Y(_4732_)
);

FILL FILL_0__15077_ (
);

AND2X2 _15362_ (
    .A(_4142__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_4318_)
);

FILL FILL360240x266760 (
);

FILL FILL187720x0 (
);

FILL FILL237880x167960 (
);

FILL FILL277400x276640 (
);

FILL FILL_1__14817_ (
);

FILL FILL290320x98800 (
);

AND2X2 _16987_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_5918_)
);

OR2X2 _16567_ (
    .A(_5504_),
    .B(_5497_),
    .Y(_5505_)
);

OR2X2 _16147_ (
    .A(_5090_),
    .B(_5089_),
    .Y(_5091_)
);

FILL FILL108680x158080 (
);

DFFSR _11282_ (
    .CLK(clk_bF$buf44),
    .D(_1389_[20]),
    .Q(\datapath_1.regfile_1.regOut[22] [20]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL_0__17643_ (
);

FILL FILL_0__17223_ (
);

AND2X2 _8489_ (
    .A(_24_),
    .B(_23_),
    .Y(_3_[10])
);

DFFSR _9850_ (
    .CLK(clk_bF$buf39),
    .D(_663_[7]),
    .Q(\datapath_1.regfile_1.regOut[11] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

OR2X2 _9430_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_530__bF$buf3),
    .Y(_512_)
);

OR2X2 _9010_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .B(_332__bF$buf3),
    .Y(_292_)
);

INVX1 _12487_ (
    .A(\control_1.reg_state.dout [1]),
    .Y(_2092_)
);

DFFSR _12067_ (
    .CLK(clk_bF$buf46),
    .D(_1785_[31]),
    .Q(\datapath_1.regfile_1.regOut[28] [31]),
    .R(rst_bF$buf97),
    .S(vdd)
);

FILL FILL_1__14150_ (
);

FILL FILL_0__18848_ (
);

OR2X2 _18713_ (
    .A(_7617_),
    .B(_7616_),
    .Y(_7618_)
);

FILL FILL_0__18428_ (
);

FILL FILL_0__13983_ (
);

FILL FILL294120x98800 (
);

FILL FILL460560x69160 (
);

FILL FILL258400x222300 (
);

FILL FILL_1__9172_ (
);

FILL FILL139840x93860 (
);

FILL FILL_1__15775_ (
);

FILL FILL_1__10070_ (
);

FILL FILL_0__14768_ (
);

OR2X2 _14633_ (
    .A(vdd),
    .B(\datapath_1.a [2]),
    .Y(_3808_)
);

OR2X2 _14213_ (
    .A(\datapath_1.Data [23]),
    .B(_3605__bF$buf4),
    .Y(_3587_)
);

FILL FILL451440x0 (
);

FILL FILL44080x39520 (
);

FILL FILL129960x276640 (
);

FILL FILL300960x9880 (
);

FILL FILL_0__18181_ (
);

AND2X2 _15838_ (
    .A(_4142__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_4787_)
);

AND2X2 _15418_ (
    .A(_4373_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd2 [2])
);

AND2X2 _10973_ (
    .A(_1300_),
    .B(_1299_),
    .Y(_1257_[21])
);

FILL FILL_1__17921_ (
);

AND2X2 _10553_ (
    .A(_1080_),
    .B(_1079_),
    .Y(_1059_[10])
);

OR2X2 _10133_ (
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .Y(_925_)
);

FILL FILL_0__16914_ (
);

AND2X2 _19251_ (
    .A(_6262__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_8148_)
);

FILL FILL117040x64220 (
);

DFFSR _8701_ (
    .CLK(clk_bF$buf81),
    .D(_69_[19]),
    .Q(\datapath_1.regfile_1.regOut[2] [19]),
    .R(rst_bF$buf19),
    .S(vdd)
);

FILL FILL_0__9067_ (
);

OR2X2 _11758_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .B(_1718__bF$buf1),
    .Y(_1704_)
);

OR2X2 _11338_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .B(_1520__bF$buf1),
    .Y(_1484_)
);

FILL FILL_1__13001_ (
);

FILL FILL_0__12834_ (
);

FILL FILL_0__12414_ (
);

OR2X2 _15591_ (
    .A(_4543_),
    .B(_4540_),
    .Y(_4544_)
);

FILL FILL28880x98800 (
);

AND2X2 _15171_ (
    .A(_4127_),
    .B(_4128_),
    .Y(_4129_)
);

FILL FILL153520x54340 (
);

OR2X2 _9906_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_749_)
);

FILL FILL_1__8863_ (
);

FILL FILL113240x177840 (
);

FILL FILL_1__14626_ (
);

FILL FILL_0__13619_ (
);

OR2X2 _13904_ (
    .A(\datapath_1.a [29]),
    .B(_3342__bF$buf2),
    .Y(_3336_)
);

FILL FILL_1__17098_ (
);

OR2X2 _16796_ (
    .A(_5729_),
    .B(_5728_),
    .Y(_5730_)
);

OR2X2 _16376_ (
    .A(_5301_),
    .B(_5316_),
    .Y(_5317_)
);

OR2X2 _11091_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_1359_)
);

FILL FILL_0__17872_ (
);

FILL FILL_0__17032_ (
);

DFFSR _12296_ (
    .CLK(clk_bF$buf56),
    .D(_1917_[2]),
    .Q(\datapath_1.regfile_1.regOut[30] [2]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL_1__19244_ (
);

OR2X2 _18942_ (
    .A(_7843_),
    .B(_7840_),
    .Y(_7844_)
);

FILL FILL_0__18237_ (
);

OR2X2 _18522_ (
    .A(_7426_),
    .B(_7429_),
    .Y(_7430_)
);

AND2X2 _18102_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_7017_)
);

FILL FILL_0__13372_ (
);

FILL FILL354160x251940 (
);

FILL FILL_0__8758_ (
);

OR2X2 _10609_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_1124__bF$buf1),
    .Y(_1118_)
);

AND2X2 _19307_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_8203_)
);

FILL FILL288800x271700 (
);

DFFSR _14862_ (
    .CLK(clk_bF$buf40),
    .D(_3870_[10]),
    .Q(_2_[10]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL_0__14577_ (
);

FILL FILL_0__14157_ (
);

OR2X2 _14442_ (
    .A(memoryOutData[24]),
    .B(_3737__bF$buf2),
    .Y(_3721_)
);

OR2X2 _14022_ (
    .A(_3438_),
    .B(_3435_),
    .Y(\datapath_1.alu_1.ALUInB [14])
);

FILL FILL279680x375440 (
);

FILL FILL363280x64220 (
);

FILL FILL411920x217360 (
);

OR2X2 _15647_ (
    .A(_4597_),
    .B(_4598_),
    .Y(_4599_)
);

OR2X2 _15227_ (
    .A(_4182_),
    .B(_4184_),
    .Y(_4185_)
);

OR2X2 _10782_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_1193_)
);

FILL FILL184680x335920 (
);

DFFSR _10362_ (
    .CLK(clk_bF$buf10),
    .D(_927_[3]),
    .Q(\datapath_1.regfile_1.regOut[15] [3]),
    .R(rst_bF$buf16),
    .S(vdd)
);

FILL FILL_0__10077_ (
);

FILL FILL_0__16723_ (
);

FILL FILL443080x232180 (
);

FILL FILL_0__19195_ (
);

AND2X2 _19480_ (
    .A(_8355_),
    .B(_8354_),
    .Y(_8320_[17])
);

FILL FILL12160x123500 (
);

AND2X2 _19060_ (
    .A(_6321__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_7960_)
);

AND2X2 _8930_ (
    .A(_258_),
    .B(_257_),
    .Y(_201_[28])
);

AND2X2 _8510_ (
    .A(_38_),
    .B(_37_),
    .Y(_3_[17])
);

FILL FILL_0__9296_ (
);

AND2X2 _11987_ (
    .A(_1816_),
    .B(_1815_),
    .Y(_1785_[15])
);

FILL FILL_1__18935_ (
);

AND2X2 _11567_ (
    .A(_1596_),
    .B(_1595_),
    .Y(_1587_[4])
);

DFFSR _11147_ (
    .CLK(clk_bF$buf21),
    .D(_1323_[14]),
    .Q(\datapath_1.regfile_1.regOut[21] [14]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL_1__13650_ (
);

FILL FILL_1__13230_ (
);

FILL FILL_0__17508_ (
);

FILL FILL_0__12223_ (
);

FILL FILL76000x54340 (
);

FILL FILL195320x207480 (
);

DFFSR _9715_ (
    .CLK(clk_bF$buf1),
    .D(_597_[1]),
    .Q(\datapath_1.regfile_1.regOut[10] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL377720x118560 (
);

FILL FILL_0__13848_ (
);

FILL FILL_0__13428_ (
);

AND2X2 _13713_ (
    .A(_3087__bF$buf2),
    .B(\datapath_1.ALUResult [17]),
    .Y(_3191_)
);

OR2X2 _16185_ (
    .A(_5128_),
    .B(_5097_),
    .Y(_5129_)
);

FILL FILL_1__9877_ (
);

FILL FILL_0__17681_ (
);

FILL FILL_0__17261_ (
);

FILL FILL354920x0 (
);

OR2X2 _14918_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [11]),
    .Y(_3958_)
);

FILL FILL487160x113620 (
);

FILL FILL_0__18886_ (
);

OR2X2 _18751_ (
    .A(_7654_),
    .B(_7655_),
    .Y(_7656_)
);

FILL FILL_0__18466_ (
);

OR2X2 _18331_ (
    .A(_7241_),
    .B(_7240_),
    .Y(_7242_)
);

FILL FILL_0__18046_ (
);

FILL FILL_0__13181_ (
);

FILL FILL_0__8987_ (
);

AND2X2 _10838_ (
    .A(_1230_),
    .B(_1229_),
    .Y(_1191_[19])
);

AND2X2 _10418_ (
    .A(_1010_),
    .B(_1009_),
    .Y(_993_[8])
);

FILL FILL388360x88920 (
);

FILL FILL343520x326040 (
);

DFFSR _19536_ (
    .CLK(clk_bF$buf38),
    .D(_8320_[13]),
    .Q(\datapath_1.regfile_1.regOut[0] [13]),
    .R(rst_bF$buf51),
    .S(vdd)
);

AND2X2 _19116_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_8015_)
);

AND2X2 _14671_ (
    .A(_3833_),
    .B(_3832_),
    .Y(_3804_[14])
);

FILL FILL_0__14386_ (
);

AND2X2 _14251_ (
    .A(_3613_),
    .B(_3612_),
    .Y(_3606_[3])
);

FILL FILL255360x291460 (
);

FILL FILL_1__16598_ (
);

FILL FILL_1__16178_ (
);

OR2X2 _15876_ (
    .A(_4822_),
    .B(_4823_),
    .Y(_4824_)
);

OR2X2 _15456_ (
    .A(_4407_),
    .B(_4410_),
    .Y(_4411_)
);

OAI21X1 _15036_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .C(_4024_),
    .Y(_4025_)
);

OR2X2 _10591_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .B(_1124__bF$buf2),
    .Y(_1106_)
);

OR2X2 _10171_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .B(_926__bF$buf2),
    .Y(_886_)
);

FILL FILL_0__16112_ (
);

FILL FILL428640x177840 (
);

FILL FILL373920x148200 (
);

FILL FILL259920x172900 (
);

DFFSR _11796_ (
    .CLK(clk_bF$buf63),
    .D(_1653_[18]),
    .Q(\datapath_1.regfile_1.regOut[26] [18]),
    .R(rst_bF$buf58),
    .S(vdd)
);

OR2X2 _11376_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_1509_)
);

FILL FILL_0__17737_ (
);

OR2X2 _17602_ (
    .A(_6509_),
    .B(_6524_),
    .Y(_6525_)
);

FILL FILL_0__17317_ (
);

FILL FILL_0__12872_ (
);

FILL FILL_0__12032_ (
);

AND2X2 _9944_ (
    .A(_774_),
    .B(_773_),
    .Y(_729_[22])
);

AND2X2 _9524_ (
    .A(_554_),
    .B(_553_),
    .Y(_531_[11])
);

AND2X2 _9104_ (
    .A(_334_),
    .B(_397_),
    .Y(_333_[0])
);

FILL FILL_1__8481_ (
);

FILL FILL_1__19109_ (
);

AND2X2 _18807_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_7711_)
);

FILL FILL_0_BUFX2_insert241 (
);

FILL FILL405840x202540 (
);

FILL FILL_0_BUFX2_insert242 (
);

FILL FILL_0_BUFX2_insert243 (
);

FILL FILL_0_BUFX2_insert244 (
);

AND2X2 _13942_ (
    .A(_3350__bF$buf1),
    .B(_2_[3]),
    .Y(_3370_)
);

FILL FILL_0_BUFX2_insert245 (
);

FILL FILL_0__13237_ (
);

OR2X2 _13522_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [11]),
    .Y(_3036_)
);

FILL FILL431680x44460 (
);

NOR2X1 _13102_ (
    .A(_2270_),
    .B(_2498_),
    .Y(_2656_)
);

FILL FILL_0_BUFX2_insert247 (
);

FILL FILL_0_BUFX2_insert249 (
);

BUFX2 BUFX2_insert1160 (
    .A(_8385_),
    .Y(_8385__bF$buf4)
);

BUFX2 BUFX2_insert1161 (
    .A(_8385_),
    .Y(_8385__bF$buf3)
);

BUFX2 BUFX2_insert1162 (
    .A(_8385_),
    .Y(_8385__bF$buf2)
);

FILL FILL_0__17490_ (
);

FILL FILL_0__17070_ (
);

BUFX2 BUFX2_insert1163 (
    .A(_8385_),
    .Y(_8385__bF$buf1)
);

BUFX2 BUFX2_insert1164 (
    .A(_8385_),
    .Y(_8385__bF$buf0)
);

BUFX2 BUFX2_insert1165 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf4 )
);

BUFX2 BUFX2_insert1166 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf3 )
);

BUFX2 BUFX2_insert1167 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf2 )
);

BUFX2 BUFX2_insert1168 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf1 )
);

BUFX2 BUFX2_insert1169 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf0 )
);

DFFSR _14727_ (
    .CLK(clk_bF$buf16),
    .D(_3804_[4]),
    .Q(\datapath_1.a [4]),
    .R(rst_bF$buf15),
    .S(vdd)
);

OR2X2 _14307_ (
    .A(\datapath_1.ALUResult [22]),
    .B(_3671__bF$buf3),
    .Y(_3651_)
);

BUFX2 BUFX2_insert980 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf0 )
);

BUFX2 BUFX2_insert981 (
    .A(_6302_),
    .Y(_6302__bF$buf4)
);

BUFX2 BUFX2_insert982 (
    .A(_6302_),
    .Y(_6302__bF$buf3)
);

BUFX2 BUFX2_insert983 (
    .A(_6302_),
    .Y(_6302__bF$buf2)
);

FILL FILL278920x158080 (
);

BUFX2 BUFX2_insert984 (
    .A(_6302_),
    .Y(_6302__bF$buf1)
);

BUFX2 BUFX2_insert985 (
    .A(_6302_),
    .Y(_6302__bF$buf0)
);

OR2X2 _17199_ (
    .A(_6123_),
    .B(_6126_),
    .Y(_6127_)
);

BUFX2 BUFX2_insert986 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf4)
);

BUFX2 BUFX2_insert987 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf3)
);

BUFX2 BUFX2_insert988 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf2)
);

BUFX2 BUFX2_insert989 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf1)
);

FILL FILL147440x266760 (
);

FILL FILL_0__18695_ (
);

OR2X2 _18980_ (
    .A(_7880_),
    .B(_7879_),
    .Y(_7881_)
);

OR2X2 _18560_ (
    .A(_7464_),
    .B(_7467_),
    .Y(_7468_)
);

OR2X2 _18140_ (
    .A(_7053_),
    .B(_7046_),
    .Y(_7054_)
);

FILL FILL_0__8796_ (
);

FILL FILL478800x59280 (
);

DFFSR _10647_ (
    .CLK(clk_bF$buf32),
    .D(_1059_[30]),
    .Q(\datapath_1.regfile_1.regOut[17] [30]),
    .R(rst_bF$buf42),
    .S(vdd)
);

OR2X2 _10227_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_923_)
);

FILL FILL_0__11723_ (
);

FILL FILL_0__11303_ (
);

FILL FILL196080x291460 (
);

AND2X2 _19345_ (
    .A(_6326__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_8241_)
);

FILL FILL187720x360620 (
);

FILL FILL_0__14195_ (
);

DFFSR _14480_ (
    .CLK(clk_bF$buf23),
    .D(_3672_[15]),
    .Q(\datapath_1.Data [15]),
    .R(rst_bF$buf33),
    .S(vdd)
);

OR2X2 _14060_ (
    .A(_3469_),
    .B(_3470_),
    .Y(_3471_)
);

FILL FILL373920x375440 (
);

FILL FILL_1__13515_ (
);

FILL FILL88920x123500 (
);

AND2X2 _15685_ (
    .A(_4151__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_4636_)
);

AND2X2 _15265_ (
    .A(_4222_),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .Y(_4223_)
);

FILL FILL300200x266760 (
);

FILL FILL19760x88920 (
);

FILL FILL_0__16761_ (
);

FILL FILL_0__16341_ (
);

FILL FILL69160x187720 (
);

OR2X2 _11185_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .B(_1454__bF$buf1),
    .Y(_1402_)
);

FILL FILL_0__17966_ (
);

FILL FILL_0__17546_ (
);

AND2X2 _17831_ (
    .A(_6282__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [7]),
    .Y(_6750_)
);

AND2X2 _17411_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_6336_)
);

FILL FILL228000x29640 (
);

FILL FILL_0__12261_ (
);

FILL FILL318440x148200 (
);

OR2X2 _9753_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_667_)
);

DFFSR _9333_ (
    .CLK(clk_bF$buf49),
    .D(_399_[6]),
    .Q(\datapath_1.regfile_1.regOut[7] [6]),
    .R(rst_bF$buf106),
    .S(vdd)
);

FILL FILL_1__19338_ (
);

AND2X2 _18616_ (
    .A(_6232__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_7523_)
);

FILL FILL_0__13886_ (
);

FILL FILL_0__13466_ (
);

OR2X2 _13751_ (
    .A(_3223_),
    .B(_3220_),
    .Y(\datapath_1.mux_pcsrc.dout [22])
);

FILL FILL_0__13046_ (
);

OR2X2 _13331_ (
    .A(_2403_),
    .B(_2400_),
    .Y(_2872_)
);

AND2X2 _14956_ (
    .A(_3983_),
    .B(_3982_),
    .Y(_3936_[23])
);

AND2X2 _14536_ (
    .A(_3763_),
    .B(_3762_),
    .Y(_3738_[12])
);

FILL FILL475000x266760 (
);

OR2X2 _14116_ (
    .A(_3517_),
    .B(_3518_),
    .Y(_3519_)
);

FILL FILL_0__15612_ (
);

FILL FILL_0__18084_ (
);

FILL FILL269800x79040 (
);

DFFSR _10876_ (
    .CLK(clk_bF$buf34),
    .D(_1191_[1]),
    .Q(\datapath_1.regfile_1.regOut[19] [1]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _10456_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_1058__bF$buf3),
    .Y(_1036_)
);

FILL FILL_1__17404_ (
);

OR2X2 _10036_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .B(_860__bF$buf4),
    .Y(_816_)
);

FILL FILL_0__11952_ (
);

FILL FILL_0__11112_ (
);

FILL FILL375440x345800 (
);

FILL FILL_0__19289_ (
);

AND2X2 _19154_ (
    .A(_6321__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_8053_)
);

OR2X2 _8604_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_81_)
);

FILL FILL289560x4940 (
);

FILL FILL_1__13744_ (
);

FILL FILL_0__12737_ (
);

INVX1 _12602_ (
    .A(_2166_),
    .Y(_2167_)
);

AND2X2 _15494_ (
    .A(_4239__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_4448_)
);

AND2X2 _15074_ (
    .A(_4060_),
    .B(_4045_),
    .Y(_4061_)
);

AND2X2 _9809_ (
    .A(_704_),
    .B(_703_),
    .Y(_663_[20])
);

FILL FILL_1__8766_ (
);

FILL FILL_0__16990_ (
);

FILL FILL501600x74100 (
);

FILL FILL_0__16570_ (
);

FILL FILL_0__16150_ (
);

FILL FILL177840x103740 (
);

FILL FILL_1__14949_ (
);

OR2X2 _13807_ (
    .A(_3271_),
    .B(_3268_),
    .Y(\datapath_1.mux_pcsrc.dout [30])
);

FILL FILL278160x311220 (
);

FILL FILL72960x153140 (
);

AND2X2 _16699_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_5634_)
);

OR2X2 _16279_ (
    .A(_5220_),
    .B(_5217_),
    .Y(_5221_)
);

FILL FILL_1__18362_ (
);

FILL FILL295640x321100 (
);

AND2X2 _17640_ (
    .A(_6229__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_6562_)
);

FILL FILL_0__17355_ (
);

FILL FILL95000x118560 (
);

OR2X2 _17220_ (
    .A(_6145_),
    .B(_6146_),
    .Y(_6147_)
);

FILL FILL_0__12070_ (
);

FILL FILL431680x187720 (
);

DFFSR _9982_ (
    .CLK(clk_bF$buf33),
    .D(_729_[10]),
    .Q(\datapath_1.regfile_1.regOut[12] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

OR2X2 _9562_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .B(_596__bF$buf4),
    .Y(_580_)
);

OR2X2 _9142_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .B(_398__bF$buf2),
    .Y(_360_)
);

FILL FILL471200x296400 (
);

OR2X2 _12199_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(_1982__bF$buf3),
    .Y(_1918_)
);

FILL FILL_0__10803_ (
);

FILL FILL277400x83980 (
);

FILL FILL116280x163020 (
);

AND2X2 _18845_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_7748_)
);

FILL FILL_0_BUFX2_insert621 (
);

OR2X2 _18425_ (
    .A(_7334_),
    .B(_7333_),
    .Y(_7335_)
);

FILL FILL_0_BUFX2_insert622 (
);

OR2X2 _18005_ (
    .A(_6920_),
    .B(_6919_),
    .Y(_6921_)
);

FILL FILL_0_BUFX2_insert623 (
);

OR2X2 _13980_ (
    .A(_3402_),
    .B(_3399_),
    .Y(\datapath_1.alu_1.ALUInB [8])
);

FILL FILL_0_BUFX2_insert624 (
);

FILL FILL_0__13695_ (
);

FILL FILL_0__13275_ (
);

AND2X2 _13560_ (
    .A(_3061_),
    .B(_3060_),
    .Y(_1_[23])
);

FILL FILL_0_BUFX2_insert625 (
);

NAND2X1 _13140_ (
    .A(_2691_),
    .B(_2689_),
    .Y(_2692_)
);

FILL FILL_0_BUFX2_insert627 (
);

FILL FILL_0_BUFX2_insert629 (
);

FILL FILL_0__19501_ (
);

FILL FILL224200x256880 (
);

FILL FILL_1__15067_ (
);

OR2X2 _14765_ (
    .A(vdd),
    .B(_2_[3]),
    .Y(_3876_)
);

DFFSR _14345_ (
    .CLK(clk_bF$buf50),
    .D(_3606_[9]),
    .Q(ALUOut[9]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL247000x340860 (
);

FILL FILL_0__15841_ (
);

FILL FILL351880x163020 (
);

AND2X2 _10685_ (
    .A(_1148_),
    .B(_1147_),
    .Y(_1125_[11])
);

AND2X2 _10265_ (
    .A(_928_),
    .B(_991_),
    .Y(_927_[0])
);

FILL FILL_0__16626_ (
);

OR2X2 _16911_ (
    .A(_5842_),
    .B(_5841_),
    .Y(_5843_)
);

FILL FILL_0__16206_ (
);

FILL FILL_0__11341_ (
);

AND2X2 _19383_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_8278_)
);

DFFSR _8833_ (
    .CLK(clk_bF$buf25),
    .D(_135_[22]),
    .Q(\datapath_1.regfile_1.regOut[3] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

BUFX2 _8413_ (
    .A(_1_[21]),
    .Y(memoryAddress[21])
);

FILL FILL144400x88920 (
);

FILL FILL_0__12966_ (
);

NAND2X1 _12831_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2396_)
);

FILL FILL_0__12546_ (
);

OR2X2 _12411_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_2039_)
);

FILL FILL103360x59280 (
);

INVX2 _9618_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .Y(_662_)
);

FILL FILL74480x123500 (
);

FILL FILL_1__14758_ (
);

AND2X2 _13616_ (
    .A(_3089__bF$buf0),
    .B(gnd),
    .Y(_3108_)
);

OR2X2 _16088_ (
    .A(_5025_),
    .B(_5032_),
    .Y(_5033_)
);

FILL FILL_1__18591_ (
);

FILL FILL_0__17584_ (
);

FILL FILL_0__17164_ (
);

FILL FILL440800x202540 (
);

FILL FILL131480x222300 (
);

FILL FILL427120x113620 (
);

AND2X2 _9791_ (
    .A(_692_),
    .B(_691_),
    .Y(_663_[14])
);

FILL FILL_1__16904_ (
);

AND2X2 _9371_ (
    .A(_472_),
    .B(_471_),
    .Y(_465_[3])
);

FILL FILL440040x108680 (
);

FILL FILL271320x103740 (
);

FILL FILL_1__19376_ (
);

FILL FILL_0__10612_ (
);

FILL FILL_1__14091_ (
);

AND2X2 _18654_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_7560_)
);

OR2X2 _18234_ (
    .A(_7143_),
    .B(_7146_),
    .Y(_7147_)
);

FILL FILL_0__19310_ (
);

FILL FILL_0__9411_ (
);

FILL FILL_1__15296_ (
);

OR2X2 _19439_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [4]),
    .Y(_8328_)
);

OR2X2 _19019_ (
    .A(_7919_),
    .B(_7918_),
    .Y(_7920_)
);

DFFSR _14994_ (
    .CLK(clk_bF$buf92),
    .D(_3936_[13]),
    .Q(\datapath_1.mux_iord.din0 [13]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL_0__14289_ (
);

OR2X2 _14574_ (
    .A(memoryOutData[25]),
    .B(_3803__bF$buf4),
    .Y(_3789_)
);

AND2X2 _14154_ (
    .A(_3547_),
    .B(_3546_),
    .Y(\datapath_1.mux_wd3.dout [3])
);

FILL FILL15960x187720 (
);

FILL FILL338960x261820 (
);

FILL FILL22040x59280 (
);

FILL FILL_0__15230_ (
);

FILL FILL351880x256880 (
);

FILL FILL186200x187720 (
);

FILL FILL_1__13609_ (
);

OR2X2 _15779_ (
    .A(_4727_),
    .B(_4728_),
    .Y(_4729_)
);

AND2X2 _15359_ (
    .A(_4225__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_4315_)
);

DFFSR _10494_ (
    .CLK(clk_bF$buf108),
    .D(_993_[6]),
    .Q(\datapath_1.regfile_1.regOut[16] [6]),
    .R(rst_bF$buf66),
    .S(vdd)
);

OR2X2 _10074_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_841_)
);

FILL FILL_0__16855_ (
);

FILL FILL_0__16435_ (
);

OR2X2 _16720_ (
    .A(_5654_),
    .B(_5651_),
    .Y(_5655_)
);

FILL FILL29640x44460 (
);

FILL FILL_0__16015_ (
);

AND2X2 _16300_ (
    .A(_4234__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_5242_)
);

FILL FILL_0__11990_ (
);

FILL FILL15200x311220 (
);

OR2X2 _19192_ (
    .A(_8089_),
    .B(_8086_),
    .Y(_8090_)
);

FILL FILL97280x217360 (
);

FILL FILL231800x330980 (
);

FILL FILL349600x133380 (
);

AND2X2 _8642_ (
    .A(_106_),
    .B(_105_),
    .Y(_69_[18])
);

FILL FILL212800x167960 (
);

AND2X2 _11699_ (
    .A(_1664_),
    .B(_1663_),
    .Y(_1653_[5])
);

FILL FILL_1__18227_ (
);

DFFSR _11279_ (
    .CLK(clk_bF$buf53),
    .D(_1389_[17]),
    .Q(\datapath_1.regfile_1.regOut[22] [17]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL505400x237120 (
);

OR2X2 _17925_ (
    .A(_6839_),
    .B(_6842_),
    .Y(_6843_)
);

OR2X2 _17505_ (
    .A(_6428_),
    .B(_6415_),
    .Y(_6429_)
);

OR2X2 _12640_ (
    .A(_2202_),
    .B(_2204_),
    .Y(_2205_)
);

FILL FILL_0__12355_ (
);

OR2X2 _12220_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .B(_1982__bF$buf1),
    .Y(_1932_)
);

FILL FILL235600x251940 (
);

DFFSR _9847_ (
    .CLK(clk_bF$buf101),
    .D(_663_[4]),
    .Q(\datapath_1.regfile_1.regOut[11] [4]),
    .R(rst_bF$buf54),
    .S(vdd)
);

OR2X2 _9427_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .B(_530__bF$buf3),
    .Y(_510_)
);

OR2X2 _9007_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .B(_332__bF$buf4),
    .Y(_290_)
);

FILL FILL285000x306280 (
);

FILL FILL180120x128440 (
);

FILL FILL_1__14567_ (
);

FILL FILL271320x330980 (
);

AND2X2 _13845_ (
    .A(_3296_),
    .B(_3295_),
    .Y(\datapath_1.alu_1.ALUInA [9])
);

OR2X2 _13425_ (
    .A(_2157__bF$buf1),
    .B(_2959_),
    .Y(_2960_)
);

AOI22X1 _13005_ (
    .A(_2320_),
    .B(_2379__bF$buf3),
    .C(_2548_),
    .D(_2318_),
    .Y(_2565_)
);

FILL FILL213560x54340 (
);

FILL FILL427880x108680 (
);

FILL FILL145920x29640 (
);

FILL FILL_0__14921_ (
);

FILL FILL_0__14501_ (
);

FILL FILL295640x0 (
);

OR2X2 _9180_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .Y(_385_)
);

FILL FILL_0__15706_ (
);

FILL FILL_0__10421_ (
);

OR2X2 _18883_ (
    .A(_7784_),
    .B(_7785_),
    .Y(_7786_)
);

FILL FILL_0__18598_ (
);

FILL FILL_0__18178_ (
);

OR2X2 _18463_ (
    .A(_7371_),
    .B(_7370_),
    .Y(_7372_)
);

AND2X2 _18043_ (
    .A(_6312__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_6959_)
);

FILL FILL424840x54340 (
);

FILL FILL217360x54340 (
);

FILL FILL_1__12633_ (
);

FILL FILL328320x153140 (
);

DFFSR _11911_ (
    .CLK(clk_bF$buf87),
    .D(_1719_[4]),
    .Q(\datapath_1.regfile_1.regOut[27] [4]),
    .R(rst_bF$buf2),
    .S(vdd)
);

FILL FILL_0__11626_ (
);

AND2X2 _19248_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_8145_)
);

AND2X2 _14383_ (
    .A(_3681_),
    .B(_3680_),
    .Y(_3672_[4])
);

FILL FILL44840x14820 (
);

FILL FILL104880x167960 (
);

AND2X2 _15588_ (
    .A(_4203__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_4541_)
);

INVX1 _15168_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_4126_)
);

FILL FILL250040x350740 (
);

FILL FILL_0__16664_ (
);

FILL FILL465120x19760 (
);

OR2X2 _8871_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_219_)
);

BUFX2 _8451_ (
    .A(_2_[27]),
    .Y(memoryWriteData[27])
);

FILL FILL45600x360620 (
);

FILL FILL_1__18876_ (
);

FILL FILL_1__18456_ (
);

OR2X2 _11088_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_1357_)
);

FILL FILL55480x306280 (
);

FILL FILL_0__17449_ (
);

OR2X2 _17734_ (
    .A(_6621_),
    .B(_6654_),
    .Y(_6655_)
);

FILL FILL_0__17029_ (
);

OR2X2 _17314_ (
    .A(_6239_),
    .B(_6237_),
    .Y(_6240_)
);

FILL FILL362520x266760 (
);

FILL FILL_0__12164_ (
);

FILL FILL359480x217360 (
);

AND2X2 _9656_ (
    .A(_622_),
    .B(_621_),
    .Y(_597_[12])
);

AND2X2 _9236_ (
    .A(_402_),
    .B(_401_),
    .Y(_399_[1])
);

FILL FILL_1__11904_ (
);

FILL FILL385320x350740 (
);

FILL FILL280440x172900 (
);

FILL FILL_1__14376_ (
);

AND2X2 _18939_ (
    .A(_6255__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_7841_)
);

AND2X2 _18519_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_7427_)
);

FILL FILL_0__13789_ (
);

AND2X2 _13654_ (
    .A(_3081__bF$buf0),
    .B(ALUOut[9]),
    .Y(_3140_)
);

OR2X2 _13234_ (
    .A(_2157__bF$buf3),
    .B(_2779_),
    .Y(_2780_)
);

FILL FILL162640x4940 (
);

FILL FILL272080x69160 (
);

FILL FILL_0__14310_ (
);

FILL FILL188480x286520 (
);

DFFSR _14859_ (
    .CLK(clk_bF$buf41),
    .D(_3870_[7]),
    .Q(_2_[7]),
    .R(rst_bF$buf63),
    .S(vdd)
);

OR2X2 _14439_ (
    .A(memoryOutData[23]),
    .B(_3737__bF$buf2),
    .Y(_3719_)
);

AND2X2 _14019_ (
    .A(_3350__bF$buf3),
    .B(_2_[14]),
    .Y(_3436_)
);

FILL FILL_0__15935_ (
);

OR2X2 _15800_ (
    .A(_4734_),
    .B(_4749_),
    .Y(_4750_)
);

FILL FILL_0__10650_ (
);

FILL FILL82840x79040 (
);

AND2X2 _18692_ (
    .A(_6287__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_7598_)
);

AND2X2 _18272_ (
    .A(_6221__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_7184_)
);

FILL FILL429400x227240 (
);

FILL FILL354920x281580 (
);

FILL FILL424080x182780 (
);

INVX2 _10779_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .Y(_1256_)
);

DFFSR _10359_ (
    .CLK(clk_bF$buf99),
    .D(_927_[0]),
    .Q(\datapath_1.regfile_1.regOut[15] [0]),
    .R(rst_bF$buf19),
    .S(vdd)
);

FILL FILL_1__12862_ (
);

FILL FILL_1__12022_ (
);

FILL FILL_0__11855_ (
);

FILL FILL_0__11435_ (
);

AND2X2 _11720_ (
    .A(_1678_),
    .B(_1677_),
    .Y(_1653_[12])
);

AND2X2 _11300_ (
    .A(_1458_),
    .B(_1457_),
    .Y(_1455_[1])
);

FILL FILL315400x345800 (
);

AND2X2 _19477_ (
    .A(_8353_),
    .B(_8352_),
    .Y(_8320_[16])
);

AND2X2 _19057_ (
    .A(_6206__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_7957_)
);

FILL FILL296400x301340 (
);

OR2X2 _14192_ (
    .A(\datapath_1.Data [16]),
    .B(_3605__bF$buf4),
    .Y(_3573_)
);

AND2X2 _8927_ (
    .A(_256_),
    .B(_255_),
    .Y(_201_[27])
);

AND2X2 _8507_ (
    .A(_36_),
    .B(_35_),
    .Y(_3_[16])
);

OR2X2 _12925_ (
    .A(_2166_),
    .B(_2489_),
    .Y(_2490_)
);

FILL FILL491720x207480 (
);

NAND2X1 _12505_ (
    .A(\control_1.reg_state.dout [1]),
    .B(\control_1.reg_state.dout [0]),
    .Y(_2102_)
);

FILL FILL_1_BUFX2_insert554 (
);

FILL FILL_1_BUFX2_insert556 (
);

FILL FILL_1_BUFX2_insert558 (
);

AND2X2 _15397_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_4353_)
);

FILL FILL_1__17480_ (
);

FILL FILL_0__16053_ (
);

OR2X2 _8680_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_134__bF$buf4),
    .Y(_132_)
);

FILL FILL111720x256880 (
);

FILL FILL235600x321100 (
);

OR2X2 _17963_ (
    .A(_6878_),
    .B(_6879_),
    .Y(_6880_)
);

FILL FILL_0__17678_ (
);

BUFX2 BUFX2_insert224 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf4 )
);

OR2X2 _17543_ (
    .A(_6464_),
    .B(_6465_),
    .Y(_6466_)
);

BUFX2 BUFX2_insert225 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf3 )
);

BUFX2 BUFX2_insert226 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf2 )
);

OR2X2 _17123_ (
    .A(_6050_),
    .B(_6051_),
    .Y(_6052_)
);

BUFX2 BUFX2_insert227 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf1 )
);

BUFX2 BUFX2_insert228 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf0 )
);

FILL FILL_0__12393_ (
);

BUFX2 BUFX2_insert229 (
    .A(_4187_),
    .Y(_4187__bF$buf4)
);

FILL FILL134520x340860 (
);

FILL FILL85880x355680 (
);

FILL FILL90440x83980 (
);

OR2X2 _9885_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_735_)
);

DFFSR _9465_ (
    .CLK(clk_bF$buf75),
    .D(_465_[9]),
    .Q(\datapath_1.regfile_1.regOut[8] [9]),
    .R(rst_bF$buf27),
    .S(vdd)
);

OR2X2 _9045_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_315_)
);

FILL FILL115520x177840 (
);

FILL FILL_1__11713_ (
);

FILL FILL_0__10706_ (
);

FILL FILL_1__14185_ (
);

OR2X2 _18748_ (
    .A(_7649_),
    .B(_7652_),
    .Y(_7653_)
);

OR2X2 _18328_ (
    .A(_7238_),
    .B(_7234_),
    .Y(_7239_)
);

OR2X2 _13883_ (
    .A(\datapath_1.a [22]),
    .B(_3342__bF$buf4),
    .Y(_3322_)
);

AND2X2 _13463_ (
    .A(_2995_),
    .B(_2835_),
    .Y(_2996_)
);

FILL FILL_0__13178_ (
);

OR2X2 _13043_ (
    .A(_2285_),
    .B(_2259_),
    .Y(_2600_)
);

FILL FILL_0__9505_ (
);

AND2X2 _14668_ (
    .A(_3831_),
    .B(_3830_),
    .Y(_3804_[13])
);

AND2X2 _14248_ (
    .A(_3611_),
    .B(_3610_),
    .Y(_3606_[2])
);

FILL FILL_0__15744_ (
);

FILL FILL_0__15324_ (
);

OR2X2 _18081_ (
    .A(_6992_),
    .B(_6995_),
    .Y(_6996_)
);

FILL FILL163400x9880 (
);

FILL FILL9120x247000 (
);

FILL FILL50920x187720 (
);

FILL FILL_1__17956_ (
);

FILL FILL301720x301340 (
);

OR2X2 _10588_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_1124__bF$buf2),
    .Y(_1104_)
);

OR2X2 _10168_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .B(_926__bF$buf4),
    .Y(_884_)
);

FILL FILL_0__16949_ (
);

FILL FILL_0__16529_ (
);

OR2X2 _16814_ (
    .A(_5747_),
    .B(_5746_),
    .Y(_5748_)
);

FILL FILL_0__11244_ (
);

FILL FILL373160x167960 (
);

OR2X2 _19286_ (
    .A(_8181_),
    .B(_8182_),
    .Y(_8183_)
);

FILL FILL460560x172900 (
);

OR2X2 _8736_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_149_)
);

FILL FILL110200x98800 (
);

FILL FILL_1__13036_ (
);

FILL FILL104880x237120 (
);

FILL FILL_0__12869_ (
);

INVX1 _12734_ (
    .A(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2299_)
);

DFFSR _12314_ (
    .CLK(clk_bF$buf44),
    .D(_1917_[20]),
    .Q(\datapath_1.regfile_1.regOut[30] [20]),
    .R(rst_bF$buf16),
    .S(vdd)
);

FILL FILL_0__12029_ (
);

FILL FILL_1__8898_ (
);

FILL FILL14440x123500 (
);

FILL FILL_0__16282_ (
);

AND2X2 _13939_ (
    .A(_3344__bF$buf2),
    .B(gnd),
    .Y(_3367_)
);

OR2X2 _13519_ (
    .A(IorD_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [10]),
    .Y(_3034_)
);

FILL FILL_1__15602_ (
);

FILL FILL449160x153140 (
);

FILL FILL504640x370500 (
);

FILL FILL320720x19760 (
);

OR2X2 _17772_ (
    .A(_6690_),
    .B(_6691_),
    .Y(_6692_)
);

FILL FILL_0__17067_ (
);

NAND3X1 _17352_ (
    .A(_6227_),
    .B(_6201_),
    .C(_6214_),
    .Y(_6278_)
);

FILL FILL354160x113620 (
);

FILL FILL113240x19760 (
);

OR2X2 _9694_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .B(_662__bF$buf0),
    .Y(_648_)
);

OR2X2 _9274_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .B(_464__bF$buf1),
    .Y(_428_)
);

FILL FILL_1__11102_ (
);

FILL FILL_0__10935_ (
);

OR2X2 _10800_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_1205_)
);

OR2X2 _18977_ (
    .A(_7874_),
    .B(_7877_),
    .Y(_7878_)
);

AND2X2 _18557_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_7465_)
);

AND2X2 _18137_ (
    .A(_6211__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_7051_)
);

AND2X2 _13692_ (
    .A(_3087__bF$buf1),
    .B(\datapath_1.ALUResult [14]),
    .Y(_3173_)
);

XOR2X1 _13272_ (
    .A(_2790_),
    .B(_2802_),
    .Y(_2816_)
);

FILL FILL_0__19213_ (
);

FILL FILL288040x360620 (
);

FILL FILL_1__12727_ (
);

FILL FILL489440x113620 (
);

FILL FILL_0__9314_ (
);

OR2X2 _14897_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [4]),
    .Y(_3944_)
);

DFFSR _14477_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[12]),
    .Q(\datapath_1.Data [12]),
    .R(rst_bF$buf85),
    .S(vdd)
);

OR2X2 _14057_ (
    .A(_3468_),
    .B(_3465_),
    .Y(\datapath_1.alu_1.ALUInB [19])
);

FILL FILL302480x79040 (
);

FILL FILL_0__15973_ (
);

FILL FILL_0__15553_ (
);

FILL FILL_0__15133_ (
);

FILL FILL328320x316160 (
);

FILL FILL415720x321100 (
);

AND2X2 _10397_ (
    .A(_996_),
    .B(_995_),
    .Y(_993_[1])
);

FILL FILL_1__17345_ (
);

FILL FILL345800x326040 (
);

FILL FILL_1__12480_ (
);

OR2X2 _16623_ (
    .A(_5559_),
    .B(_5556_),
    .Y(_5560_)
);

AND2X2 _16203_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [15]),
    .Y(_5146_)
);

FILL FILL_0__11473_ (
);

FILL FILL_0__11053_ (
);

FILL FILL340480x281580 (
);

OR2X2 _19095_ (
    .A(_7994_),
    .B(_7991_),
    .Y(_7995_)
);

DFFSR _8965_ (
    .CLK(clk_bF$buf43),
    .D(_201_[25]),
    .Q(\datapath_1.regfile_1.regOut[4] [25]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL257640x291460 (
);

OR2X2 _8545_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .B(_68__bF$buf4),
    .Y(_62_)
);

FILL FILL_1__13685_ (
);

OR2X2 _17828_ (
    .A(_6743_),
    .B(_6746_),
    .Y(_6747_)
);

OR2X2 _17408_ (
    .A(_6283_),
    .B(_6333_),
    .Y(_6334_)
);

OR2X2 _12963_ (
    .A(_2523_),
    .B(_2525_),
    .Y(_2526_)
);

FILL FILL_0__12678_ (
);

FILL FILL_1_BUFX2_insert933 (
);

INVX1 _12543_ (
    .A(\control_1.op [1]),
    .Y(_2132_)
);

OR2X2 _12123_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_1887_)
);

FILL FILL_1_BUFX2_insert935 (
);

FILL FILL_1_BUFX2_insert937 (
);

FILL FILL380000x256880 (
);

FILL FILL_0__18904_ (
);

FILL FILL77520x311220 (
);

AND2X2 _13748_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [22]),
    .Y(_3221_)
);

AOI22X1 _13328_ (
    .A(_2868_),
    .B(_2379__bF$buf2),
    .C(_2593_),
    .D(_2411_),
    .Y(_2869_)
);

FILL FILL17480x64220 (
);

FILL FILL_0__14824_ (
);

FILL FILL436240x345800 (
);

BUFX2 BUFX2_insert600 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf39)
);

FILL FILL94240x227240 (
);

BUFX2 BUFX2_insert601 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf38)
);

BUFX2 BUFX2_insert602 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf37)
);

BUFX2 BUFX2_insert603 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf36)
);

BUFX2 BUFX2_insert604 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf35)
);

OR2X2 _17581_ (
    .A(_6503_),
    .B(_6501_),
    .Y(_6504_)
);

FILL FILL_0__17296_ (
);

BUFX2 BUFX2_insert605 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf34)
);

OR2X2 _17161_ (
    .A(_6088_),
    .B(_6081_),
    .Y(_6089_)
);

BUFX2 BUFX2_insert606 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf33)
);

BUFX2 BUFX2_insert607 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf32)
);

BUFX2 BUFX2_insert608 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf31)
);

BUFX2 BUFX2_insert609 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf30)
);

FILL FILL145920x158080 (
);

FILL FILL221160x321100 (
);

DFFSR _9083_ (
    .CLK(clk_bF$buf37),
    .D(_267_[14]),
    .Q(\datapath_1.regfile_1.regOut[5] [14]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_0__15609_ (
);

FILL FILL_0__10744_ (
);

FILL FILL_0__10324_ (
);

AND2X2 _18786_ (
    .A(_6229__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_7690_)
);

OR2X2 _18366_ (
    .A(_7269_),
    .B(_7276_),
    .Y(_7277_)
);

OR2X2 _13081_ (
    .A(_2635_),
    .B(_2615_),
    .Y(_2636_)
);

FILL FILL206720x64220 (
);

FILL FILL_0__19442_ (
);

FILL FILL238640x103740 (
);

FILL FILL310840x370500 (
);

FILL FILL337440x83980 (
);

FILL FILL_0__9543_ (
);

OR2X2 _11814_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_1721_)
);

FILL FILL_0__9123_ (
);

FILL FILL98040x335920 (
);

OR2X2 _14286_ (
    .A(\datapath_1.ALUResult [15]),
    .B(_3671__bF$buf2),
    .Y(_3637_)
);

FILL FILL72200x281580 (
);

FILL FILL_0__15782_ (
);

FILL FILL376200x192660 (
);

FILL FILL286520x326040 (
);

FILL FILL434720x14820 (
);

FILL FILL_1__17994_ (
);

FILL FILL_1__17574_ (
);

FILL FILL478040x59280 (
);

FILL FILL253840x187720 (
);

FILL FILL_0__16567_ (
);

AND2X2 _16852_ (
    .A(_4187__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_5785_)
);

AND2X2 _16432_ (
    .A(_4142__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_5372_)
);

FILL FILL_0__16147_ (
);

OR2X2 _16012_ (
    .A(_4957_),
    .B(_4956_),
    .Y(_4958_)
);

FILL FILL272080x256880 (
);

FILL FILL_1__9704_ (
);

FILL FILL137560x49400 (
);

AND2X2 _8774_ (
    .A(_174_),
    .B(_173_),
    .Y(_135_[19])
);

FILL FILL30400x143260 (
);

FILL FILL_1__10602_ (
);

FILL FILL411920x88920 (
);

FILL FILL_1__13074_ (
);

AND2X2 _17637_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_6559_)
);

OR2X2 _17217_ (
    .A(_6140_),
    .B(_6143_),
    .Y(_6144_)
);

OR2X2 _12772_ (
    .A(_2326_),
    .B(_2336_),
    .Y(_2337_)
);

FILL FILL_0__12487_ (
);

OR2X2 _12352_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .B(_2048__bF$buf3),
    .Y(_2000_)
);

FILL FILL_0__18713_ (
);

DFFSR _9979_ (
    .CLK(clk_bF$buf39),
    .D(_729_[7]),
    .Q(\datapath_1.regfile_1.regOut[12] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

OR2X2 _9559_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_596__bF$buf1),
    .Y(_578_)
);

OR2X2 _9139_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .B(_398__bF$buf2),
    .Y(_358_)
);

FILL FILL_1__14699_ (
);

FILL FILL222680x9880 (
);

FILL FILL_0_BUFX2_insert590 (
);

FILL FILL_0_BUFX2_insert592 (
);

AND2X2 _13977_ (
    .A(_3350__bF$buf1),
    .B(_2_[8]),
    .Y(_3400_)
);

FILL FILL_0_BUFX2_insert594 (
);

AND2X2 _13557_ (
    .A(_3059_),
    .B(_3058_),
    .Y(_1_[22])
);

AOI21X1 _13137_ (
    .A(_2288_),
    .B(_2504_),
    .C(_2688_),
    .Y(_2689_)
);

FILL FILL_0_BUFX2_insert596 (
);

FILL FILL_0_BUFX2_insert597 (
);

FILL FILL_0_BUFX2_insert598 (
);

FILL FILL_0_BUFX2_insert599 (
);

FILL FILL348080x242060 (
);

FILL FILL_0__14633_ (
);

AND2X2 _17390_ (
    .A(_6315__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_6316_)
);

FILL FILL180120x34580 (
);

FILL FILL_1__16425_ (
);

FILL FILL_1__11560_ (
);

FILL FILL_0__15418_ (
);

OR2X2 _15703_ (
    .A(_4653_),
    .B(_4650_),
    .Y(_4654_)
);

FILL FILL_0__10553_ (
);

FILL FILL_0__10133_ (
);

OR2X2 _18595_ (
    .A(_7501_),
    .B(_7494_),
    .Y(_7502_)
);

FILL FILL251560x370500 (
);

AND2X2 _18175_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_7089_)
);

FILL FILL452960x123500 (
);

FILL FILL260680x9880 (
);

FILL FILL391400x251940 (
);

OR2X2 _16908_ (
    .A(_5838_),
    .B(_5839_),
    .Y(_5840_)
);

FILL FILL_0__11758_ (
);

OR2X2 _11623_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_1652__bF$buf3),
    .Y(_1634_)
);

OR2X2 _11203_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .B(_1454__bF$buf0),
    .Y(_1414_)
);

FILL FILL4560x138320 (
);

FILL FILL125400x182780 (
);

OR2X2 _14095_ (
    .A(_3499_),
    .B(_3500_),
    .Y(_3501_)
);

FILL FILL243960x4940 (
);

FILL FILL289560x14820 (
);

FILL FILL222680x133380 (
);

FILL FILL_0__15171_ (
);

FILL FILL69160x370500 (
);

XNOR2X1 _12828_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2393_)
);

OR2X2 _12408_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_2037_)
);

FILL FILL82080x365560 (
);

FILL FILL505400x123500 (
);

FILL FILL377720x345800 (
);

FILL FILL401280x321100 (
);

FILL FILL_0__16796_ (
);

AND2X2 _16661_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_5597_)
);

FILL FILL_0__16376_ (
);

AND2X2 _16241_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [15]),
    .Y(_5184_)
);

FILL FILL_0__11091_ (
);

FILL FILL_1__9513_ (
);

FILL FILL266760x88920 (
);

FILL FILL450680x88920 (
);

DFFSR _8583_ (
    .CLK(clk_bF$buf32),
    .D(_3_[30]),
    .Q(\datapath_1.regfile_1.regOut[1] [30]),
    .R(rst_bF$buf93),
    .S(vdd)
);

FILL FILL43320x182780 (
);

FILL FILL_1__10411_ (
);

AND2X2 _17866_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_6784_)
);

AND2X2 _17446_ (
    .A(_6328__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_6371_)
);

AND2X2 _17026_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_5956_)
);

OR2X2 _12581_ (
    .A(vdd),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2151_)
);

AND2X2 _12161_ (
    .A(_1912_),
    .B(_1911_),
    .Y(_1851_[30])
);

FILL FILL480320x83980 (
);

FILL FILL_0__18942_ (
);

AND2X2 _9788_ (
    .A(_690_),
    .B(_689_),
    .Y(_663_[13])
);

AND2X2 _9368_ (
    .A(_470_),
    .B(_469_),
    .Y(_465_[2])
);

FILL FILL_0__10609_ (
);

FILL FILL380760x311220 (
);

OR2X2 _13786_ (
    .A(_3253_),
    .B(_3250_),
    .Y(\datapath_1.mux_pcsrc.dout [27])
);

AND2X2 _13366_ (
    .A(_2904_),
    .B(_2892_),
    .Y(_2905_)
);

FILL FILL370120x271700 (
);

FILL FILL29640x276640 (
);

FILL FILL_0__19307_ (
);

CLKBUF1 CLKBUF1_insert1170 (
    .A(clk),
    .Y(clk_hier0_bF$buf9)
);

FILL FILL456000x286520 (
);

CLKBUF1 CLKBUF1_insert1171 (
    .A(clk),
    .Y(clk_hier0_bF$buf8)
);

CLKBUF1 CLKBUF1_insert1172 (
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

FILL FILL_0__14442_ (
);

CLKBUF1 CLKBUF1_insert1173 (
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

FILL FILL_0__14022_ (
);

CLKBUF1 CLKBUF1_insert1174 (
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1175 (
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1176 (
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1177 (
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1178 (
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert1179 (
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert140 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf83)
);

CLKBUF1 CLKBUF1_insert141 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf82)
);

CLKBUF1 CLKBUF1_insert142 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf81)
);

CLKBUF1 CLKBUF1_insert143 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf80)
);

FILL FILL_0__9828_ (
);

CLKBUF1 CLKBUF1_insert144 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf79)
);

FILL FILL_0__9408_ (
);

CLKBUF1 CLKBUF1_insert145 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf78)
);

CLKBUF1 CLKBUF1_insert146 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf77)
);

CLKBUF1 CLKBUF1_insert147 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf76)
);

CLKBUF1 CLKBUF1_insert148 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf75)
);

CLKBUF1 CLKBUF1_insert149 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf74)
);

FILL FILL118560x163020 (
);

AND2X2 _15932_ (
    .A(_4142__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_4879_)
);

FILL FILL_0__15647_ (
);

OR2X2 _15512_ (
    .A(_4465_),
    .B(_4458_),
    .Y(_4466_)
);

FILL FILL101080x247000 (
);

FILL FILL_0__10782_ (
);

FILL FILL_0__19480_ (
);

FILL FILL_0__19060_ (
);

FILL FILL_1__17439_ (
);

FILL FILL414200x148200 (
);

FILL FILL_1__12154_ (
);

FILL FILL32680x242060 (
);

AND2X2 _16717_ (
    .A(_4167__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_5652_)
);

FILL FILL_0__11987_ (
);

FILL FILL_0__9581_ (
);

FILL FILL_0__11567_ (
);

AND2X2 _11852_ (
    .A(_1746_),
    .B(_1745_),
    .Y(_1719_[13])
);

AND2X2 _11432_ (
    .A(_1526_),
    .B(_1525_),
    .Y(_1521_[2])
);

FILL FILL505400x350740 (
);

DFFSR _11012_ (
    .CLK(clk_bF$buf84),
    .D(_1257_[8]),
    .Q(\datapath_1.regfile_1.regOut[20] [8]),
    .R(rst_bF$buf47),
    .S(vdd)
);

AND2X2 _19189_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_8087_)
);

AND2X2 _8639_ (
    .A(_104_),
    .B(_103_),
    .Y(_69_[17])
);

FILL FILL122360x59280 (
);

FILL FILL180880x143260 (
);

XOR2X1 _12637_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2202_)
);

OR2X2 _12217_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .B(_1982__bF$buf1),
    .Y(_1930_)
);

FILL FILL289560x242060 (
);

FILL FILL_0__13713_ (
);

FILL FILL272080x326040 (
);

AND2X2 _16890_ (
    .A(_5822_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd2 [25])
);

FILL FILL_0__16185_ (
);

OR2X2 _16470_ (
    .A(_5408_),
    .B(_5407_),
    .Y(_5409_)
);

OR2X2 _16050_ (
    .A(_4995_),
    .B(_4994_),
    .Y(_4996_)
);

FILL FILL448400x167960 (
);

FILL FILL344280x365560 (
);

BUFX2 _8392_ (
    .A(_1_[0]),
    .Y(memoryAddress[0])
);

FILL FILL_0__14918_ (
);

FILL FILL_1__18397_ (
);

FILL FILL376960x113620 (
);

AND2X2 _17675_ (
    .A(_6315__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_6596_)
);

OR2X2 _17255_ (
    .A(_6178_),
    .B(_6181_),
    .Y(_6182_)
);

OR2X2 _12390_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_2025_)
);

FILL FILL_0__18331_ (
);

FILL FILL250800x153140 (
);

DFFSR _9597_ (
    .CLK(clk_bF$buf102),
    .D(_531_[12]),
    .Q(\datapath_1.regfile_1.regOut[9] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

OR2X2 _9177_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_383_)
);

FILL FILL_1__11845_ (
);

FILL FILL_0__8432_ (
);

FILL FILL_0__10838_ (
);

FILL FILL_0__10418_ (
);

AND2X2 _10703_ (
    .A(_1160_),
    .B(_1159_),
    .Y(_1125_[17])
);

FILL FILL_0_BUFX2_insert970 (
);

FILL FILL_0_BUFX2_insert972 (
);

FILL FILL_0_BUFX2_insert974 (
);

AND2X2 _13595_ (
    .A(_3089__bF$buf0),
    .B(gnd),
    .Y(_3090_)
);

OR2X2 _13175_ (
    .A(_2387__bF$buf0),
    .B(_2724_),
    .Y(_2725_)
);

FILL FILL_0_BUFX2_insert976 (
);

FILL FILL_0_BUFX2_insert977 (
);

FILL FILL_0_BUFX2_insert978 (
);

FILL FILL_0_BUFX2_insert979 (
);

OR2X2 _19401_ (
    .A(_8294_),
    .B(_8295_),
    .Y(_8296_)
);

FILL FILL373160x98800 (
);

FILL FILL_0__14671_ (
);

FILL FILL133760x222300 (
);

FILL FILL_0__9637_ (
);

FILL FILL429400x113620 (
);

DFFSR _11908_ (
    .CLK(clk_bF$buf34),
    .D(_1719_[1]),
    .Q(\datapath_1.regfile_1.regOut[27] [1]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_1__16463_ (
);

FILL FILL_1__16043_ (
);

FILL FILL68400x153140 (
);

OR2X2 _15741_ (
    .A(_4690_),
    .B(_4689_),
    .Y(_4691_)
);

FILL FILL_0__15036_ (
);

OR2X2 _15321_ (
    .A(_4277_),
    .B(_4262_),
    .Y(_4278_)
);

FILL FILL_0__10171_ (
);

FILL FILL440800x276640 (
);

FILL FILL184680x59280 (
);

OR2X2 _16946_ (
    .A(_5876_),
    .B(_5877_),
    .Y(_5878_)
);

AND2X2 _16526_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_5464_)
);

AND2X2 _16106_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_5051_)
);

DFFSR _11661_ (
    .CLK(clk_bF$buf102),
    .D(_1587_[12]),
    .Q(\datapath_1.regfile_1.regOut[25] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

FILL FILL_0__11376_ (
);

OR2X2 _11241_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_1439_)
);

FILL FILL_0__17602_ (
);

OR2X2 _8868_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_217_)
);

BUFX2 _8448_ (
    .A(_2_[24]),
    .Y(memoryWriteData[24])
);

FILL FILL_1__13168_ (
);

NOR2X1 _12866_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2431_)
);

DFFSR _12446_ (
    .CLK(clk_bF$buf87),
    .D(_1983_[23]),
    .Q(\datapath_1.regfile_1.regOut[31] [23]),
    .R(rst_bF$buf2),
    .S(vdd)
);

AND2X2 _12026_ (
    .A(_1842_),
    .B(_1841_),
    .Y(_1785_[28])
);

FILL FILL_0__18807_ (
);

FILL FILL_0__13942_ (
);

FILL FILL_0__13522_ (
);

FILL FILL_0__13102_ (
);

FILL FILL319960x24700 (
);

FILL FILL_0__8908_ (
);

FILL FILL_1__9131_ (
);

AND2X2 _17484_ (
    .A(_6328__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_6408_)
);

OR2X2 _17064_ (
    .A(_5993_),
    .B(_5986_),
    .Y(_5994_)
);

FILL FILL338200x138320 (
);

FILL FILL_0__18980_ (
);

FILL FILL_0__18560_ (
);

FILL FILL383040x242060 (
);

FILL FILL_1__16939_ (
);

OR2X2 _10932_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_1273_)
);

DFFSR _10512_ (
    .CLK(clk_bF$buf97),
    .D(_993_[24]),
    .Q(\datapath_1.regfile_1.regOut[16] [24]),
    .R(rst_bF$buf84),
    .S(vdd)
);

OR2X2 _18689_ (
    .A(_7594_),
    .B(_7593_),
    .Y(_7595_)
);

OR2X2 _18269_ (
    .A(_7177_),
    .B(_7180_),
    .Y(_7181_)
);

FILL FILL_0__19345_ (
);

OR2X2 _19210_ (
    .A(_8100_),
    .B(_8107_),
    .Y(_8108_)
);

FILL FILL146680x261820 (
);

FILL FILL_0__14060_ (
);

FILL FILL_0__9446_ (
);

FILL FILL196080x316160 (
);

AND2X2 _11717_ (
    .A(_1676_),
    .B(_1675_),
    .Y(_1653_[11])
);

FILL FILL_0__9026_ (
);

FILL FILL283480x321100 (
);

OR2X2 _14189_ (
    .A(\datapath_1.Data [15]),
    .B(_3605__bF$buf3),
    .Y(_3571_)
);

FILL FILL_1__16692_ (
);

FILL FILL63840x14820 (
);

AND2X2 _15970_ (
    .A(_4183__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_4917_)
);

FILL FILL_0__15685_ (
);

FILL FILL_0__15265_ (
);

AND2X2 _15550_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_4503_)
);

AND2X2 _15130_ (
    .A(_4029_),
    .B(_4105_),
    .Y(\datapath_1.regfile_1.regEn [14])
);

FILL FILL155800x83980 (
);

FILL FILL40280x14820 (
);

FILL FILL43320x79040 (
);

FILL FILL294880x256880 (
);

AND2X2 _16755_ (
    .A(_4239__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_5690_)
);

OR2X2 _16335_ (
    .A(_5275_),
    .B(_5274_),
    .Y(_5276_)
);

OR2X2 _11890_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .B(_1784__bF$buf4),
    .Y(_1772_)
);

OR2X2 _11470_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .B(_1586__bF$buf1),
    .Y(_1552_)
);

FILL FILL_0__11185_ (
);

OR2X2 _11050_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .B(_1388__bF$buf2),
    .Y(_1332_)
);

FILL FILL95760x247000 (
);

FILL FILL_0__17831_ (
);

FILL FILL_0__17411_ (
);

OR2X2 _8677_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .B(_134__bF$buf3),
    .Y(_130_)
);

FILL FILL129200x266760 (
);

FILL FILL298680x177840 (
);

FILL FILL67640x14820 (
);

FILL FILL266000x326040 (
);

OR2X2 _12675_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(_2239_),
    .Y(_2240_)
);

FILL FILL_1__19203_ (
);

OR2X2 _12255_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_1955_)
);

OR2X2 _18901_ (
    .A(_7796_),
    .B(_7803_),
    .Y(_7804_)
);

FILL FILL252320x350740 (
);

FILL FILL_0__13751_ (
);

FILL FILL_0__8717_ (
);

FILL FILL332120x4940 (
);

FILL FILL434720x261820 (
);

FILL FILL_1__15543_ (
);

AND2X2 _14821_ (
    .A(_3913_),
    .B(_3912_),
    .Y(_3870_[21])
);

FILL FILL_0__14116_ (
);

AND2X2 _14401_ (
    .A(_3693_),
    .B(_3692_),
    .Y(_3672_[10])
);

FILL FILL364800x266760 (
);

AND2X2 _17293_ (
    .A(_6218_),
    .B(\datapath_1.PCJump [25]),
    .Y(_6219_)
);

FILL FILL351120x4940 (
);

FILL FILL387600x350740 (
);

FILL FILL234840x74100 (
);

FILL FILL_1__11463_ (
);

OR2X2 _15606_ (
    .A(_4555_),
    .B(_4558_),
    .Y(_4559_)
);

FILL FILL_0__8890_ (
);

FILL FILL_0__10456_ (
);

OR2X2 _10741_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .B(_1190__bF$buf4),
    .Y(_1186_)
);

OR2X2 _10321_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_992__bF$buf2),
    .Y(_966_)
);

AND2X2 _18498_ (
    .A(_6272__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_7407_)
);

AND2X2 _18078_ (
    .A(_6216__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_6993_)
);

FILL FILL_0__19154_ (
);

FILL FILL350360x0 (
);

FILL FILL121600x375440 (
);

FILL FILL_1__12668_ (
);

FILL FILL118560x326040 (
);

FILL FILL_0__9255_ (
);

OR2X2 _11946_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_1789_)
);

DFFSR _11526_ (
    .CLK(clk_bF$buf29),
    .D(_1521_[6]),
    .Q(\datapath_1.regfile_1.regOut[24] [6]),
    .R(rst_bF$buf40),
    .S(vdd)
);

OR2X2 _11106_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_1369_)
);

FILL FILL104880x350740 (
);

FILL FILL278920x24700 (
);

FILL FILL_0__12602_ (
);

FILL FILL345800x212420 (
);

FILL FILL_0__15494_ (
);

FILL FILL231040x370500 (
);

FILL FILL426360x182780 (
);

FILL FILL_0__13807_ (
);

FILL FILL443840x192660 (
);

FILL FILL_0__16699_ (
);

OR2X2 _16984_ (
    .A(_5914_),
    .B(_5907_),
    .Y(_5915_)
);

AND2X2 _16564_ (
    .A(_4130__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_5502_)
);

OR2X2 _16144_ (
    .A(_5087_),
    .B(_5084_),
    .Y(_5088_)
);

FILL FILL408880x355680 (
);

FILL FILL_1__9416_ (
);

FILL FILL343520x286520 (
);

AND2X2 _8486_ (
    .A(_22_),
    .B(_21_),
    .Y(_3_[9])
);

FILL FILL_1__10734_ (
);

FILL FILL184680x227240 (
);

OR2X2 _17769_ (
    .A(_6687_),
    .B(_6688_),
    .Y(_6689_)
);

NAND3X1 _17349_ (
    .A(_6227_),
    .B(\datapath_1.PCJump [24]),
    .C(_6225_),
    .Y(_6275_)
);

AND2X2 _12484_ (
    .A(_2075_),
    .B(ALUOp[1]),
    .Y(_2076_)
);

DFFSR _12064_ (
    .CLK(clk_bF$buf74),
    .D(_1785_[28]),
    .Q(\datapath_1.regfile_1.regOut[28] [28]),
    .R(rst_bF$buf47),
    .S(vdd)
);

FILL FILL_0__18845_ (
);

AND2X2 _18710_ (
    .A(_7615_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd1 [20])
);

FILL FILL_0__18425_ (
);

FILL FILL_0__18005_ (
);

FILL FILL_0__13560_ (
);

FILL FILL_0__13140_ (
);

FILL FILL_0__8526_ (
);

AND2X2 _13689_ (
    .A(_3081__bF$buf0),
    .B(ALUOut[14]),
    .Y(_3170_)
);

NOR2X1 _13269_ (
    .A(_2644_),
    .B(_2810_),
    .Y(_2813_)
);

OR2X2 _14630_ (
    .A(vdd),
    .B(\datapath_1.a [1]),
    .Y(_3806_)
);

OR2X2 _14210_ (
    .A(\datapath_1.Data [22]),
    .B(_3605__bF$buf2),
    .Y(_3585_)
);

FILL FILL199120x54340 (
);

FILL FILL136800x340860 (
);

FILL FILL152000x24700 (
);

FILL FILL_1__16557_ (
);

AND2X2 _15835_ (
    .A(_4158__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_4784_)
);

OR2X2 _15415_ (
    .A(_4363_),
    .B(_4370_),
    .Y(_4371_)
);

AND2X2 _10970_ (
    .A(_1298_),
    .B(_1297_),
    .Y(_1257_[20])
);

FILL FILL_0__10685_ (
);

AND2X2 _10550_ (
    .A(_1078_),
    .B(_1077_),
    .Y(_1059_[9])
);

FILL FILL_0__10265_ (
);

DFFSR _10130_ (
    .CLK(clk_bF$buf88),
    .D(_795_[29]),
    .Q(\datapath_1.regfile_1.regOut[13] [29]),
    .R(rst_bF$buf112),
    .S(vdd)
);

FILL FILL240920x261820 (
);

FILL FILL277400x321100 (
);

FILL FILL_0__19383_ (
);

FILL FILL_1__18703_ (
);

OR2X2 _11755_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .B(_1718__bF$buf4),
    .Y(_1702_)
);

OR2X2 _11335_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .B(_1520__bF$buf1),
    .Y(_1482_)
);

FILL FILL_0__12831_ (
);

FILL FILL35720x177840 (
);

FILL FILL80560x281580 (
);

FILL FILL206720x158080 (
);

OR2X2 _9903_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_747_)
);

FILL FILL495520x311220 (
);

FILL FILL58520x261820 (
);

FILL FILL71440x256880 (
);

FILL FILL294880x98800 (
);

OR2X2 _13901_ (
    .A(\datapath_1.a [28]),
    .B(_3342__bF$buf4),
    .Y(_3334_)
);

FILL FILL_0__13616_ (
);

FILL FILL462840x172900 (
);

FILL FILL193800x74100 (
);

OR2X2 _16793_ (
    .A(_5726_),
    .B(_5711_),
    .Y(_5727_)
);

FILL FILL_0__16088_ (
);

OR2X2 _16373_ (
    .A(_5312_),
    .B(_5313_),
    .Y(_5314_)
);

FILL FILL427880x335920 (
);

FILL FILL12920x202540 (
);

FILL FILL205960x0 (
);

FILL FILL_1__15408_ (
);

FILL FILL115520x69160 (
);

FILL FILL_1__10543_ (
);

BUFX2 BUFX2_insert570 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf69)
);

BUFX2 BUFX2_insert571 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf68)
);

BUFX2 BUFX2_insert572 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf67)
);

BUFX2 BUFX2_insert573 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf66)
);

BUFX2 BUFX2_insert574 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf65)
);

OR2X2 _17998_ (
    .A(_6912_),
    .B(_6913_),
    .Y(_6914_)
);

AND2X2 _17578_ (
    .A(_6289__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_6501_)
);

BUFX2 BUFX2_insert575 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf64)
);

BUFX2 BUFX2_insert576 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf63)
);

AND2X2 _17158_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_6086_)
);

BUFX2 BUFX2_insert577 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf62)
);

BUFX2 BUFX2_insert578 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf61)
);

BUFX2 BUFX2_insert579 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf60)
);

FILL FILL447640x232180 (
);

AND2X2 _12293_ (
    .A(_1980_),
    .B(_1979_),
    .Y(_1917_[31])
);

FILL FILL_0__18654_ (
);

FILL FILL132240x276640 (
);

FILL FILL_1__11748_ (
);

OR2X2 _10606_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .B(_1124__bF$buf2),
    .Y(_1116_)
);

FILL FILL10640x54340 (
);

FILL FILL_0_BUFX2_insert90 (
);

FILL FILL_0_BUFX2_insert92 (
);

FILL FILL253840x0 (
);

FILL FILL_0_BUFX2_insert94 (
);

FILL FILL197600x74100 (
);

FILL FILL_0_BUFX2_insert95 (
);

FILL FILL_0_BUFX2_insert96 (
);

FILL FILL_0_BUFX2_insert97 (
);

OR2X2 _13498_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [3]),
    .Y(_3020_)
);

FILL FILL411160x44460 (
);

AND2X2 _13078_ (
    .A(_2633_),
    .B(_2625_),
    .Y(_2634_)
);

FILL FILL_0_BUFX2_insert98 (
);

FILL FILL_0_BUFX2_insert99 (
);

FILL FILL_1__15581_ (
);

FILL FILL_1__15161_ (
);

FILL FILL_0__19019_ (
);

AND2X2 _19304_ (
    .A(_6300__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_8200_)
);

FILL FILL_0__14574_ (
);

FILL FILL_0__14154_ (
);

FILL FILL_0__15779_ (
);

FILL FILL_0__15359_ (
);

OR2X2 _15644_ (
    .A(_4595_),
    .B(_4594_),
    .Y(_4596_)
);

AND2X2 _15224_ (
    .A(_4181__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_4182_)
);

FILL FILL_0__10074_ (
);

FILL FILL_0__16720_ (
);

FILL FILL_0__16300_ (
);

FILL FILL468160x256880 (
);

AND2X2 _16849_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_5782_)
);

AND2X2 _16429_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_5369_)
);

OR2X2 _16009_ (
    .A(_4954_),
    .B(_4947_),
    .Y(_4955_)
);

AND2X2 _11984_ (
    .A(_1814_),
    .B(_1813_),
    .Y(_1785_[14])
);

FILL FILL_0__9293_ (
);

FILL FILL_0__11699_ (
);

AND2X2 _11564_ (
    .A(_1594_),
    .B(_1593_),
    .Y(_1587_[3])
);

FILL FILL505400x83980 (
);

DFFSR _11144_ (
    .CLK(clk_bF$buf45),
    .D(_1323_[11]),
    .Q(\datapath_1.regfile_1.regOut[21] [11]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL_0__17925_ (
);

FILL FILL_0__12640_ (
);

FILL FILL50920x44460 (
);

OR2X2 _9712_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_662__bF$buf2),
    .Y(_660_)
);

NAND2X1 _12769_ (
    .A(_2332_),
    .B(_2333_),
    .Y(_2334_)
);

OR2X2 _12349_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .B(_2048__bF$buf1),
    .Y(_1998_)
);

AND2X2 _13710_ (
    .A(_3081__bF$buf2),
    .B(ALUOut[17]),
    .Y(_3188_)
);

FILL FILL_0__13005_ (
);

FILL FILL342760x281580 (
);

FILL FILL261440x217360 (
);

OR2X2 _16182_ (
    .A(_5122_),
    .B(_5125_),
    .Y(_5126_)
);

FILL FILL178600x227240 (
);

FILL FILL242440x375440 (
);

OR2X2 _14915_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [10]),
    .Y(_3956_)
);

AND2X2 _17387_ (
    .A(_6312__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_6313_)
);

FILL FILL246240x296400 (
);

FILL FILL_0__18463_ (
);

FILL FILL_0__18043_ (
);

FILL FILL225720x64220 (
);

FILL FILL_0__8984_ (
);

AND2X2 _10835_ (
    .A(_1228_),
    .B(_1227_),
    .Y(_1191_[18])
);

AND2X2 _10415_ (
    .A(_1008_),
    .B(_1007_),
    .Y(_993_[7])
);

FILL FILL_0__19248_ (
);

DFFSR _19533_ (
    .CLK(clk_bF$buf88),
    .D(_8320_[10]),
    .Q(\datapath_1.regfile_1.regOut[0] [10]),
    .R(rst_bF$buf37),
    .S(vdd)
);

OR2X2 _19113_ (
    .A(_8011_),
    .B(_8010_),
    .Y(_8012_)
);

FILL FILL_0__14383_ (
);

FILL FILL_0__9769_ (
);

OR2X2 _15873_ (
    .A(_4820_),
    .B(_4817_),
    .Y(_4821_)
);

FILL FILL_0__15588_ (
);

AND2X2 _15453_ (
    .A(_4142__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_4408_)
);

FILL FILL_0__15168_ (
);

FILL FILL96520x69160 (
);

NAND3X1 _15033_ (
    .A(_4018_),
    .B(_4005_),
    .C(\datapath_1.a3 [2]),
    .Y(_4022_)
);

FILL FILL229520x64220 (
);

FILL FILL_1__14908_ (
);

FILL FILL475000x158080 (
);

AND2X2 _16658_ (
    .A(_4177__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_5594_)
);

OR2X2 _16238_ (
    .A(_5179_),
    .B(_5180_),
    .Y(_5181_)
);

FILL FILL461320x182780 (
);

FILL FILL_1__18741_ (
);

DFFSR _11793_ (
    .CLK(clk_bF$buf90),
    .D(_1653_[15]),
    .Q(\datapath_1.regfile_1.regOut[26] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL_1__18321_ (
);

OR2X2 _11373_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [26]),
    .Y(_1507_)
);

FILL FILL380000x118560 (
);

FILL FILL458280x133380 (
);

FILL FILL_0__17314_ (
);

FILL FILL288800x326040 (
);

FILL FILL40280x340860 (
);

AND2X2 _9941_ (
    .A(_772_),
    .B(_771_),
    .Y(_729_[21])
);

AND2X2 _9521_ (
    .A(_552_),
    .B(_551_),
    .Y(_531_[10])
);

OR2X2 _9101_ (
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .Y(_397_)
);

XOR2X1 _12998_ (
    .A(_2325_),
    .B(_2558_),
    .Y(_2559_)
);

OR2X2 _12578_ (
    .A(vdd),
    .B(\control_1.reg_state.dout [2]),
    .Y(_2149_)
);

AND2X2 _12158_ (
    .A(_1910_),
    .B(_1909_),
    .Y(_1851_[29])
);

FILL FILL_1__14661_ (
);

FILL FILL_0__18939_ (
);

OR2X2 _18804_ (
    .A(_7707_),
    .B(_7699_),
    .Y(_7708_)
);

FILL FILL_0__18519_ (
);

FILL FILL367840x49400 (
);

FILL FILL_0__13654_ (
);

FILL FILL_0__13234_ (
);

FILL FILL75240x247000 (
);

FILL FILL398240x321100 (
);

FILL FILL_1__9263_ (
);

BUFX2 BUFX2_insert1130 (
    .A(_3350_),
    .Y(_3350__bF$buf4)
);

FILL FILL348080x172900 (
);

BUFX2 BUFX2_insert1131 (
    .A(_3350_),
    .Y(_3350__bF$buf3)
);

BUFX2 BUFX2_insert1132 (
    .A(_3350_),
    .Y(_3350__bF$buf2)
);

BUFX2 BUFX2_insert1133 (
    .A(_3350_),
    .Y(_3350__bF$buf1)
);

BUFX2 BUFX2_insert1134 (
    .A(_3350_),
    .Y(_3350__bF$buf0)
);

BUFX2 BUFX2_insert1135 (
    .A(_4135_),
    .Y(_4135__bF$buf4)
);

BUFX2 BUFX2_insert1136 (
    .A(_4135_),
    .Y(_4135__bF$buf3)
);

BUFX2 BUFX2_insert1137 (
    .A(_4135_),
    .Y(_4135__bF$buf2)
);

BUFX2 BUFX2_insert1138 (
    .A(_4135_),
    .Y(_4135__bF$buf1)
);

FILL FILL_1__15026_ (
);

BUFX2 BUFX2_insert1139 (
    .A(_4135_),
    .Y(_4135__bF$buf0)
);

DFFSR _14724_ (
    .CLK(clk_bF$buf4),
    .D(_3804_[1]),
    .Q(\datapath_1.a [1]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _14304_ (
    .A(\datapath_1.ALUResult [21]),
    .B(_3671__bF$buf1),
    .Y(_3649_)
);

BUFX2 BUFX2_insert950 (
    .A(_4065_),
    .Y(_4065__bF$buf5)
);

BUFX2 BUFX2_insert951 (
    .A(_4065_),
    .Y(_4065__bF$buf4)
);

BUFX2 BUFX2_insert952 (
    .A(_4065_),
    .Y(_4065__bF$buf3)
);

BUFX2 BUFX2_insert953 (
    .A(_4065_),
    .Y(_4065__bF$buf2)
);

BUFX2 BUFX2_insert954 (
    .A(_4065_),
    .Y(_4065__bF$buf1)
);

BUFX2 BUFX2_insert955 (
    .A(_4065_),
    .Y(_4065__bF$buf0)
);

BUFX2 BUFX2_insert956 (
    .A(_6211_),
    .Y(_6211__bF$buf4)
);

AND2X2 _17196_ (
    .A(_4228__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_6124_)
);

BUFX2 BUFX2_insert957 (
    .A(_6211_),
    .Y(_6211__bF$buf3)
);

FILL FILL_0__15800_ (
);

BUFX2 BUFX2_insert958 (
    .A(_6211_),
    .Y(_6211__bF$buf2)
);

BUFX2 BUFX2_insert959 (
    .A(_6211_),
    .Y(_6211__bF$buf1)
);

FILL FILL302480x113620 (
);

FILL FILL_0__18272_ (
);

FILL FILL450680x9880 (
);

OR2X2 _15929_ (
    .A(_4845_),
    .B(_4876_),
    .Y(_4877_)
);

AND2X2 _15509_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_4463_)
);

DFFSR _10644_ (
    .CLK(clk_bF$buf39),
    .D(_1059_[27]),
    .Q(\datapath_1.regfile_1.regOut[17] [27]),
    .R(rst_bF$buf69),
    .S(vdd)
);

OR2X2 _10224_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_921_)
);

FILL FILL_0__11720_ (
);

FILL FILL496280x167960 (
);

FILL FILL_0__11300_ (
);

AND2X2 _19342_ (
    .A(_6302__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_8238_)
);

FILL FILL_0__14192_ (
);

FILL FILL433960x4940 (
);

FILL FILL492480x14820 (
);

FILL FILL_0__9578_ (
);

FILL FILL_0__9158_ (
);

AND2X2 _11849_ (
    .A(_1744_),
    .B(_1743_),
    .Y(_1719_[12])
);

AND2X2 _11429_ (
    .A(_1524_),
    .B(_1523_),
    .Y(_1521_[1])
);

DFFSR _11009_ (
    .CLK(clk_bF$buf104),
    .D(_1257_[5]),
    .Q(\datapath_1.regfile_1.regOut[20] [5]),
    .R(rst_bF$buf25),
    .S(vdd)
);

FILL FILL_1__13932_ (
);

FILL FILL_0__12925_ (
);

FILL FILL_0__12505_ (
);

FILL FILL253840x370500 (
);

AND2X2 _15682_ (
    .A(_4203__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_4633_)
);

OR2X2 _15262_ (
    .A(_4212_),
    .B(_4219_),
    .Y(_4220_)
);

FILL FILL452960x4940 (
);

FILL FILL_1__8534_ (
);

FILL FILL76000x251940 (
);

FILL FILL11400x163020 (
);

FILL FILL6840x138320 (
);

OR2X2 _16887_ (
    .A(_5812_),
    .B(_5819_),
    .Y(_5820_)
);

OR2X2 _16467_ (
    .A(_5405_),
    .B(_5404_),
    .Y(_5406_)
);

OR2X2 _16047_ (
    .A(_4992_),
    .B(_4989_),
    .Y(_4993_)
);

FILL FILL_1__18970_ (
);

OR2X2 _11182_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .B(_1454__bF$buf1),
    .Y(_1400_)
);

FILL FILL_0__17963_ (
);

FILL FILL_0__17543_ (
);

FILL FILL_0__17123_ (
);

FILL FILL503120x108680 (
);

OR2X2 _9750_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_665_)
);

DFFSR _9330_ (
    .CLK(clk_bF$buf95),
    .D(_399_[3]),
    .Q(\datapath_1.regfile_1.regOut[7] [3]),
    .R(rst_bF$buf9),
    .S(vdd)
);

OR2X2 _12387_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_2023_)
);

FILL FILL_1__14050_ (
);

FILL FILL316160x316160 (
);

FILL FILL_0__18748_ (
);

AND2X2 _18613_ (
    .A(_6272__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_7520_)
);

FILL FILL_0__18328_ (
);

FILL FILL403560x321100 (
);

FILL FILL_0__13883_ (
);

FILL FILL_0__13043_ (
);

FILL FILL302480x340860 (
);

FILL FILL_0__8849_ (
);

FILL FILL_0__8429_ (
);

FILL FILL234080x222300 (
);

FILL FILL_1__15675_ (
);

FILL FILL_0__14668_ (
);

AND2X2 _14953_ (
    .A(_3981_),
    .B(_3980_),
    .Y(_3936_[22])
);

FILL FILL_0__14248_ (
);

AND2X2 _14533_ (
    .A(_3761_),
    .B(_3760_),
    .Y(_3738_[11])
);

OR2X2 _14113_ (
    .A(_3516_),
    .B(_3513_),
    .Y(\datapath_1.alu_1.ALUInB [27])
);

FILL FILL505400x197600 (
);

FILL FILL486400x153140 (
);

FILL FILL_1__11595_ (
);

AND2X2 _15738_ (
    .A(_4688_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd2 [7])
);

OR2X2 _15318_ (
    .A(_4274_),
    .B(_4273_),
    .Y(_4275_)
);

OR2X2 _10873_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .B(_1256__bF$buf3),
    .Y(_1254_)
);

FILL FILL_0__10588_ (
);

FILL FILL_1__17821_ (
);

OR2X2 _10453_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .B(_1058__bF$buf1),
    .Y(_1034_)
);

FILL FILL468920x326040 (
);

OR2X2 _10033_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_860__bF$buf2),
    .Y(_814_)
);

FILL FILL300200x311220 (
);

FILL FILL_0__16814_ (
);

FILL FILL_0__19286_ (
);

AND2X2 _19151_ (
    .A(_6297__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_8050_)
);

OR2X2 _8601_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_79_)
);

FILL FILL228760x29640 (
);

FILL FILL_0__9387_ (
);

DFFSR _11658_ (
    .CLK(clk_bF$buf103),
    .D(_1587_[9]),
    .Q(\datapath_1.regfile_1.regOut[25] [9]),
    .R(rst_bF$buf45),
    .S(vdd)
);

OR2X2 _11238_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_1437_)
);

FILL FILL142120x281580 (
);

FILL FILL103360x247000 (
);

FILL FILL_0__12734_ (
);

AND2X2 _15491_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_4445_)
);

AND2X2 _15071_ (
    .A(_4058_),
    .B(_4029_),
    .Y(\datapath_1.regfile_1.regEn [2])
);

FILL FILL367080x296400 (
);

FILL FILL17480x232180 (
);

AND2X2 _9806_ (
    .A(_702_),
    .B(_701_),
    .Y(_663_[19])
);

FILL FILL243200x128440 (
);

AND2X2 _13804_ (
    .A(_3087__bF$buf1),
    .B(\datapath_1.ALUResult [30]),
    .Y(_3269_)
);

FILL FILL_0__13519_ (
);

FILL FILL101840x14820 (
);

FILL FILL226480x103740 (
);

FILL FILL315400x167960 (
);

OR2X2 _16696_ (
    .A(_5616_),
    .B(_5631_),
    .Y(_5632_)
);

FILL FILL338960x153140 (
);

AND2X2 _16276_ (
    .A(_4175__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_5218_)
);

FILL FILL_1__9548_ (
);

FILL FILL_0__17772_ (
);

FILL FILL_1__10866_ (
);

FILL FILL60040x281580 (
);

FILL FILL364040x192660 (
);

DFFSR _12196_ (
    .CLK(clk_bF$buf83),
    .D(_1851_[31]),
    .Q(\datapath_1.regfile_1.regOut[29] [31]),
    .R(rst_bF$buf23),
    .S(vdd)
);

FILL FILL_1__19144_ (
);

FILL FILL_0__18977_ (
);

FILL FILL416480x360620 (
);

AND2X2 _18842_ (
    .A(_6216__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_7745_)
);

FILL FILL_0__18137_ (
);

OR2X2 _18422_ (
    .A(_7328_),
    .B(_7331_),
    .Y(_7332_)
);

OR2X2 _18002_ (
    .A(_6914_),
    .B(_6917_),
    .Y(_6918_)
);

FILL FILL_0__13692_ (
);

FILL FILL_0__13272_ (
);

FILL FILL346560x365560 (
);

FILL FILL_0__8658_ (
);

FILL FILL105640x14820 (
);

OR2X2 _10929_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_1271_)
);

DFFSR _10509_ (
    .CLK(clk_bF$buf47),
    .D(_993_[21]),
    .Q(\datapath_1.regfile_1.regOut[16] [21]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL125400x29640 (
);

AND2X2 _19207_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_8105_)
);

OR2X2 _14762_ (
    .A(vdd),
    .B(_2_[2]),
    .Y(_3874_)
);

FILL FILL_0__14057_ (
);

DFFSR _14342_ (
    .CLK(clk_bF$buf62),
    .D(_3606_[6]),
    .Q(ALUOut[6]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL421800x158080 (
);

FILL FILL72960x276640 (
);

FILL FILL78280x350740 (
);

OR2X2 _15967_ (
    .A(_4913_),
    .B(_4912_),
    .Y(_4914_)
);

AND2X2 _15547_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_4500_)
);

AND2X2 _15127_ (
    .A(_4029_),
    .B(_4103_),
    .Y(\datapath_1.regfile_1.regEn [13])
);

FILL FILL_0__10397_ (
);

AND2X2 _10682_ (
    .A(_1146_),
    .B(_1145_),
    .Y(_1125_[10])
);

FILL FILL_1__17210_ (
);

OR2X2 _10262_ (
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .Y(_991_)
);

FILL FILL_0__16623_ (
);

OR2X2 _19380_ (
    .A(_8272_),
    .B(_8274_),
    .Y(_8275_)
);

FILL FILL_0__19095_ (
);

DFFSR _8830_ (
    .CLK(clk_bF$buf81),
    .D(_135_[19]),
    .Q(\datapath_1.regfile_1.regOut[3] [19]),
    .R(rst_bF$buf101),
    .S(vdd)
);

BUFX2 _8410_ (
    .A(_1_[18]),
    .Y(memoryAddress[18])
);

FILL FILL129200x29640 (
);

FILL FILL_1__18835_ (
);

OR2X2 _11887_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .B(_1784__bF$buf3),
    .Y(_1770_)
);

OR2X2 _11467_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .B(_1586__bF$buf0),
    .Y(_1550_)
);

OR2X2 _11047_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_1388__bF$buf2),
    .Y(_1330_)
);

FILL FILL_1__13550_ (
);

FILL FILL80560x34580 (
);

FILL FILL_0__17828_ (
);

FILL FILL_0__17408_ (
);

FILL FILL440800x44460 (
);

FILL FILL_0__12123_ (
);

DFFSR _9615_ (
    .CLK(clk_bF$buf7),
    .D(_531_[30]),
    .Q(\datapath_1.regfile_1.regOut[9] [30]),
    .R(rst_bF$buf48),
    .S(vdd)
);

FILL FILL233320x44460 (
);

FILL FILL_0__13748_ (
);

FILL FILL408120x54340 (
);

FILL FILL_0__13328_ (
);

AND2X2 _13613_ (
    .A(_3084__bF$buf0),
    .B(\aluControl_1.inst [1]),
    .Y(_3105_)
);

FILL FILL160360x29640 (
);

AND2X2 _16085_ (
    .A(_4135__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_5030_)
);

FILL FILL_0__17581_ (
);

FILL FILL_0__17161_ (
);

FILL FILL_1__10675_ (
);

AND2X2 _14818_ (
    .A(_3911_),
    .B(_3910_),
    .Y(_3870_[20])
);

FILL FILL108680x98800 (
);

FILL FILL_0__18786_ (
);

OR2X2 _18651_ (
    .A(_7555_),
    .B(_7556_),
    .Y(_7557_)
);

FILL FILL_0__18366_ (
);

AND2X2 _18231_ (
    .A(_6236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_7144_)
);

FILL FILL371640x29640 (
);

FILL FILL_0__13081_ (
);

FILL FILL_0__8467_ (
);

OR2X2 _10738_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .B(_1190__bF$buf1),
    .Y(_1184_)
);

FILL FILL164160x29640 (
);

OR2X2 _10318_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_992__bF$buf1),
    .Y(_964_)
);

FILL FILL_0__11814_ (
);

OR2X2 _19436_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_8326_)
);

INVX1 _19016_ (
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_7917_)
);

DFFSR _14991_ (
    .CLK(clk_bF$buf92),
    .D(_3936_[10]),
    .Q(\datapath_1.mux_iord.din0 [10]),
    .R(rst_bF$buf29),
    .S(vdd)
);

OR2X2 _14571_ (
    .A(memoryOutData[24]),
    .B(_3803__bF$buf4),
    .Y(_3787_)
);

AND2X2 _14151_ (
    .A(_3545_),
    .B(_3544_),
    .Y(\datapath_1.mux_wd3.dout [2])
);

FILL FILL385320x242060 (
);

FILL FILL446120x212420 (
);

FILL FILL42560x64220 (
);

FILL FILL_1__16498_ (
);

OR2X2 _15776_ (
    .A(_4722_),
    .B(_4725_),
    .Y(_4726_)
);

AND2X2 _15356_ (
    .A(_4160__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_4312_)
);

DFFSR _10491_ (
    .CLK(clk_bF$buf56),
    .D(_993_[3]),
    .Q(\datapath_1.regfile_1.regOut[16] [3]),
    .R(rst_bF$buf49),
    .S(vdd)
);

OR2X2 _10071_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_839_)
);

FILL FILL_1__8628_ (
);

FILL FILL151240x83980 (
);

FILL FILL_0__16432_ (
);

FILL FILL_0__16012_ (
);

FILL FILL148960x261820 (
);

FILL FILL252320x197600 (
);

FILL FILL326040x93860 (
);

FILL FILL85120x118560 (
);

AND2X2 _11696_ (
    .A(_1662_),
    .B(_1661_),
    .Y(_1653_[4])
);

FILL FILL_1__18644_ (
);

DFFSR _11276_ (
    .CLK(clk_bF$buf85),
    .D(_1389_[14]),
    .Q(\datapath_1.regfile_1.regOut[22] [14]),
    .R(rst_bF$buf109),
    .S(vdd)
);

AND2X2 _17922_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_6840_)
);

FILL FILL_0__17637_ (
);

FILL FILL_0__17217_ (
);

OR2X2 _17502_ (
    .A(_6425_),
    .B(_6424_),
    .Y(_6426_)
);

FILL FILL_0__12772_ (
);

FILL FILL63080x14820 (
);

DFFSR _9844_ (
    .CLK(clk_bF$buf93),
    .D(_663_[1]),
    .Q(\datapath_1.regfile_1.regOut[11] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

OR2X2 _9424_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .B(_530__bF$buf0),
    .Y(_508_)
);

OR2X2 _9004_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .B(_332__bF$buf2),
    .Y(_288_)
);

FILL FILL_1__19009_ (
);

FILL FILL66120x79040 (
);

FILL FILL315400x237120 (
);

FILL FILL155040x83980 (
);

OR2X2 _18707_ (
    .A(_7597_),
    .B(_7612_),
    .Y(_7613_)
);

FILL FILL_0__13977_ (
);

AND2X2 _13842_ (
    .A(_3294_),
    .B(_3293_),
    .Y(\datapath_1.alu_1.ALUInA [8])
);

FILL FILL_0__13557_ (
);

XOR2X1 _13422_ (
    .A(_2390_),
    .B(_2852_),
    .Y(_2957_)
);

XOR2X1 _13002_ (
    .A(_2321_),
    .B(_2542_),
    .Y(_2562_)
);

FILL FILL237880x242060 (
);

FILL FILL63840x88920 (
);

FILL FILL15200x247000 (
);

FILL FILL351120x316160 (
);

FILL FILL_0__17390_ (
);

FILL FILL_1__15349_ (
);

FILL FILL_1__10484_ (
);

INVX2 _14627_ (
    .A(vdd),
    .Y(_3869_)
);

FILL FILL253840x74100 (
);

OR2X2 _14207_ (
    .A(\datapath_1.Data [21]),
    .B(_3605__bF$buf4),
    .Y(_3583_)
);

AND2X2 _17099_ (
    .A(_4183__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_6028_)
);

FILL FILL_1__19182_ (
);

FILL FILL230280x74100 (
);

OR2X2 _18880_ (
    .A(_7781_),
    .B(_7782_),
    .Y(_7783_)
);

FILL FILL_0__18595_ (
);

OR2X2 _18460_ (
    .A(_7368_),
    .B(_7367_),
    .Y(_7369_)
);

OR2X2 _18040_ (
    .A(_6955_),
    .B(_6948_),
    .Y(_6956_)
);

FILL FILL280440x291460 (
);

FILL FILL165680x4940 (
);

AND2X2 _10967_ (
    .A(_1296_),
    .B(_1295_),
    .Y(_1257_[19])
);

AND2X2 _10547_ (
    .A(_1076_),
    .B(_1075_),
    .Y(_1059_[8])
);

DFFSR _10127_ (
    .CLK(clk_bF$buf75),
    .D(_795_[26]),
    .Q(\datapath_1.regfile_1.regOut[13] [26]),
    .R(rst_bF$buf27),
    .S(vdd)
);

FILL FILL_1__12210_ (
);

FILL FILL_0__16908_ (
);

FILL FILL_0__11203_ (
);

OR2X2 _19245_ (
    .A(_8134_),
    .B(_8141_),
    .Y(_8142_)
);

FILL FILL472720x340860 (
);

FILL FILL_0__14095_ (
);

AND2X2 _14380_ (
    .A(_3679_),
    .B(_3678_),
    .Y(_3672_[3])
);

FILL FILL453720x177840 (
);

FILL FILL389880x158080 (
);

FILL FILL_1__13415_ (
);

FILL FILL_0__12408_ (
);

AND2X2 _15585_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_4538_)
);

AND2X2 _15165_ (
    .A(_4004_),
    .B(_4043_),
    .Y(\datapath_1.regfile_1.regEn [29])
);

FILL FILL275880x276640 (
);

FILL FILL_0__16661_ (
);

FILL FILL_0__16241_ (
);

OR2X2 _11085_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_1355_)
);

FILL FILL_0__17866_ (
);

FILL FILL_0__17446_ (
);

OR2X2 _17731_ (
    .A(_6651_),
    .B(_6644_),
    .Y(_6652_)
);

AND2X2 _17311_ (
    .A(_6236__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_6237_)
);

FILL FILL278160x24700 (
);

FILL FILL233320x370500 (
);

FILL FILL347320x118560 (
);

AND2X2 _9653_ (
    .A(_620_),
    .B(_619_),
    .Y(_597_[11])
);

AND2X2 _9233_ (
    .A(_400_),
    .B(_463_),
    .Y(_399_[0])
);

FILL FILL_1__14793_ (
);

AND2X2 _18936_ (
    .A(_6259__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_7838_)
);

AND2X2 _18516_ (
    .A(_6206__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_7424_)
);

FILL FILL41800x375440 (
);

FILL FILL_0__13366_ (
);

AND2X2 _13651_ (
    .A(_3089__bF$buf1),
    .B(gnd),
    .Y(_3138_)
);

AND2X2 _13231_ (
    .A(_2777_),
    .B(_2767_),
    .Y(_2778_)
);

FILL FILL256880x222300 (
);

FILL FILL345800x286520 (
);

FILL FILL_1__9395_ (
);

FILL FILL255360x98800 (
);

FILL FILL_1__15998_ (
);

FILL FILL_1__10293_ (
);

DFFSR _14856_ (
    .CLK(clk_bF$buf38),
    .D(_3870_[4]),
    .Q(_2_[4]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _14436_ (
    .A(memoryOutData[22]),
    .B(_3737__bF$buf4),
    .Y(_3717_)
);

AND2X2 _14016_ (
    .A(_3344__bF$buf0),
    .B(gnd),
    .Y(_3433_)
);

FILL FILL_0_CLKBUF1_insert200 (
);

FILL FILL_0_CLKBUF1_insert202 (
);

FILL FILL_0__15512_ (
);

FILL FILL_0_CLKBUF1_insert204 (
);

FILL FILL_0_CLKBUF1_insert205 (
);

FILL FILL_0_CLKBUF1_insert206 (
);

FILL FILL_0_CLKBUF1_insert207 (
);

FILL FILL_0_CLKBUF1_insert208 (
);

FILL FILL_0_CLKBUF1_insert209 (
);

FILL FILL3800x335920 (
);

DFFSR _10776_ (
    .CLK(clk_bF$buf109),
    .D(_1125_[30]),
    .Q(\datapath_1.regfile_1.regOut[18] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

OR2X2 _10356_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_989_)
);

FILL FILL_1__17304_ (
);

FILL FILL465880x19760 (
);

FILL FILL_0__11432_ (
);

FILL FILL_0__19189_ (
);

AND2X2 _19474_ (
    .A(_8351_),
    .B(_8350_),
    .Y(_8320_[15])
);

AND2X2 _19054_ (
    .A(_6236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_7954_)
);

AND2X2 _8924_ (
    .A(_254_),
    .B(_253_),
    .Y(_201_[26])
);

AND2X2 _8504_ (
    .A(_34_),
    .B(_33_),
    .Y(_3_[15])
);

FILL FILL_1__18509_ (
);

FILL FILL186960x9880 (
);

FILL FILL_1_BUFX2_insert521 (
);

NOR2X1 _12922_ (
    .A(_2355_),
    .B(_2357_),
    .Y(_2487_)
);

FILL FILL_0__12637_ (
);

FILL FILL_0__12217_ (
);

NOR3X1 _12502_ (
    .A(_2099_),
    .B(\control_1.reg_state.dout [1]),
    .C(\control_1.reg_state.dout [0]),
    .Y(PCWrite)
);

FILL FILL_1_BUFX2_insert529 (
);

AND2X2 _15394_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_4350_)
);

OR2X2 _9709_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .B(_662__bF$buf4),
    .Y(_658_)
);

FILL FILL_0__16890_ (
);

FILL FILL_0__16470_ (
);

FILL FILL_0__16050_ (
);

FILL FILL_1__14429_ (
);

AND2X2 _13707_ (
    .A(_3089__bF$buf2),
    .B(gnd),
    .Y(_3186_)
);

FILL FILL149720x4940 (
);

OR2X2 _16599_ (
    .A(_5532_),
    .B(_5535_),
    .Y(_5536_)
);

AND2X2 _16179_ (
    .A(_4239__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_5123_)
);

FILL FILL_1__18262_ (
);

FILL FILL288040x118560 (
);

FILL FILL375440x123500 (
);

AND2X2 _17960_ (
    .A(_6282__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [9]),
    .Y(_6877_)
);

FILL FILL_0__17255_ (
);

AND2X2 _17540_ (
    .A(_6463_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd1 [2])
);

FILL FILL82840x281580 (
);

OR2X2 _17120_ (
    .A(_6048_),
    .B(_6045_),
    .Y(_6049_)
);

OR2X2 _9882_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_733_)
);

DFFSR _9462_ (
    .CLK(clk_bF$buf104),
    .D(_465_[6]),
    .Q(\datapath_1.regfile_1.regOut[8] [6]),
    .R(rst_bF$buf8),
    .S(vdd)
);

OR2X2 _9042_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_313_)
);

FILL FILL73720x256880 (
);

OR2X2 _12099_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_1871_)
);

FILL FILL_0__10703_ (
);

AND2X2 _18745_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_7650_)
);

INVX1 _18325_ (
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_7236_)
);

OR2X2 _13880_ (
    .A(\datapath_1.a [21]),
    .B(_3342__bF$buf4),
    .Y(_3320_)
);

FILL FILL_0__13595_ (
);

FILL FILL_0__13175_ (
);

AND2X2 _13460_ (
    .A(_2992_),
    .B(_2727_),
    .Y(_2993_)
);

AND2X2 _13040_ (
    .A(_2597_),
    .B(_2595_),
    .Y(_2598_)
);

FILL FILL200640x350740 (
);

FILL FILL_0__19401_ (
);

FILL FILL193040x74100 (
);

FILL FILL_1__12915_ (
);

FILL FILL_0__9922_ (
);

FILL FILL199880x266760 (
);

FILL FILL127680x306280 (
);

AND2X2 _14665_ (
    .A(_3829_),
    .B(_3828_),
    .Y(_3804_[12])
);

AND2X2 _14245_ (
    .A(_3609_),
    .B(_3608_),
    .Y(_3606_[1])
);

FILL FILL_0__15741_ (
);

FILL FILL380760x133380 (
);

OR2X2 _10585_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .B(_1124__bF$buf0),
    .Y(_1102_)
);

OR2X2 _10165_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_926__bF$buf3),
    .Y(_882_)
);

FILL FILL_0__16946_ (
);

OR2X2 _16811_ (
    .A(_5744_),
    .B(_5743_),
    .Y(_5745_)
);

FILL FILL_0__16106_ (
);

OR2X2 _19283_ (
    .A(_8179_),
    .B(_8176_),
    .Y(_8180_)
);

OR2X2 _8733_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_147_)
);

FILL FILL_0__12866_ (
);

INVX1 _12731_ (
    .A(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2296_)
);

FILL FILL_0__12026_ (
);

DFFSR _12311_ (
    .CLK(clk_bF$buf6),
    .D(_1917_[17]),
    .Q(\datapath_1.regfile_1.regOut[30] [17]),
    .R(rst_bF$buf6),
    .S(vdd)
);

AND2X2 _9938_ (
    .A(_770_),
    .B(_769_),
    .Y(_729_[20])
);

AND2X2 _9518_ (
    .A(_550_),
    .B(_549_),
    .Y(_531_[9])
);

FILL FILL_1__14238_ (
);

AND2X2 _13936_ (
    .A(_3352__bF$buf1),
    .B(\aluControl_1.inst [0]),
    .Y(_3365_)
);

OR2X2 _13516_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [9]),
    .Y(_3032_)
);

FILL FILL310840x128440 (
);

FILL FILL_0__17484_ (
);

FILL FILL_1__10578_ (
);

FILL FILL88160x172900 (
);

FILL FILL10640x138320 (
);

FILL FILL333640x212420 (
);

OR2X2 _9691_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .B(_662__bF$buf4),
    .Y(_646_)
);

FILL FILL_1__16804_ (
);

OR2X2 _9271_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .B(_464__bF$buf1),
    .Y(_426_)
);

FILL FILL_1__19276_ (
);

FILL FILL27360x281580 (
);

FILL FILL_0__18689_ (
);

AND2X2 _18974_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_7875_)
);

FILL FILL263720x217360 (
);

AND2X2 _18554_ (
    .A(_6302__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_7462_)
);

FILL FILL_0__18269_ (
);

AND2X2 _18134_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_7048_)
);

FILL FILL_0__19210_ (
);

FILL FILL_0__11717_ (
);

OR2X2 _19339_ (
    .A(_8234_),
    .B(_8233_),
    .Y(_8235_)
);

OR2X2 _14894_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [3]),
    .Y(_3942_)
);

FILL FILL_0__14189_ (
);

DFFSR _14474_ (
    .CLK(clk_bF$buf2),
    .D(_3672_[9]),
    .Q(\datapath_1.Data [9]),
    .R(rst_bF$buf33),
    .S(vdd)
);

AND2X2 _14054_ (
    .A(_3350__bF$buf4),
    .B(_2_[19]),
    .Y(_3466_)
);

FILL FILL110960x98800 (
);

FILL FILL_0__15550_ (
);

FILL FILL_0__15130_ (
);

FILL FILL354160x370500 (
);

FILL FILL382280x103740 (
);

FILL FILL299440x113620 (
);

FILL FILL140600x93860 (
);

AND2X2 _15679_ (
    .A(_4172__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_4630_)
);

AND2X2 _15259_ (
    .A(_4216_),
    .B(_4144_),
    .Y(_4217_)
);

FILL FILL449160x276640 (
);

FILL FILL_1__17762_ (
);

AND2X2 _10394_ (
    .A(_994_),
    .B(_1057_),
    .Y(_993_[0])
);

FILL FILL98800x227240 (
);

FILL FILL_0__16755_ (
);

AND2X2 _16620_ (
    .A(_4187__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_5557_)
);

FILL FILL_0__16335_ (
);

OR2X2 _16200_ (
    .A(_5142_),
    .B(_5139_),
    .Y(_5143_)
);

FILL FILL_0__11890_ (
);

FILL FILL_0__11470_ (
);

FILL FILL101840x256880 (
);

AND2X2 _19092_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_7992_)
);

DFFSR _8962_ (
    .CLK(clk_bF$buf91),
    .D(_201_[22]),
    .Q(\datapath_1.regfile_1.regOut[4] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

OR2X2 _8542_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_68__bF$buf0),
    .Y(_60_)
);

OR2X2 _11599_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_1652__bF$buf1),
    .Y(_1618_)
);

FILL FILL459800x64220 (
);

FILL FILL_1__18127_ (
);

OR2X2 _11179_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .B(_1454__bF$buf3),
    .Y(_1398_)
);

FILL FILL297160x187720 (
);

AND2X2 _17825_ (
    .A(_6321__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_6744_)
);

FILL FILL155800x326040 (
);

OR2X2 _17405_ (
    .A(_6325_),
    .B(_6330_),
    .Y(_6331_)
);

FILL FILL_1_BUFX2_insert901 (
);

AND2X2 _12960_ (
    .A(_2521_),
    .B(_2522_),
    .Y(_2523_)
);

FILL FILL_0__12675_ (
);

FILL FILL105640x177840 (
);

FILL FILL_0__12255_ (
);

OR2X2 _12540_ (
    .A(_2122_),
    .B(_2128_),
    .Y(_2129_)
);

OR2X2 _12120_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_1885_)
);

FILL FILL269040x14820 (
);

FILL FILL_0__18901_ (
);

FILL FILL_1_BUFX2_insert909 (
);

INVX2 _9747_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .Y(_728_)
);

DFFSR _9327_ (
    .CLK(clk_bF$buf99),
    .D(_399_[0]),
    .Q(\datapath_1.regfile_1.regOut[7] [0]),
    .R(rst_bF$buf72),
    .S(vdd)
);

FILL FILL144400x93860 (
);

FILL FILL437000x0 (
);

AND2X2 _13745_ (
    .A(_3081__bF$buf2),
    .B(ALUOut[22]),
    .Y(_3218_)
);

INVX1 _13325_ (
    .A(_2411_),
    .Y(_2866_)
);

FILL FILL_0__14821_ (
);

FILL FILL443080x217360 (
);

FILL FILL_0__14401_ (
);

FILL FILL_1__9489_ (
);

FILL FILL412680x59280 (
);

DFFSR _9080_ (
    .CLK(clk_bF$buf71),
    .D(_267_[11]),
    .Q(\datapath_1.regfile_1.regOut[5] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL_0__15606_ (
);

FILL FILL_0__10741_ (
);

FILL FILL276640x256880 (
);

AND2X2 _18783_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_7687_)
);

FILL FILL_0__18078_ (
);

AND2X2 _18363_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_7274_)
);

FILL FILL367080x49400 (
);

FILL FILL_0__8599_ (
);

FILL FILL_1__12113_ (
);

FILL FILL_0__9960_ (
);

FILL FILL_0__11946_ (
);

FILL FILL_0__9540_ (
);

INVX2 _11811_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .Y(_1784_)
);

FILL FILL_0__11106_ (
);

NOR2X1 _19148_ (
    .A(_6310__bF$buf4),
    .B(_8046_),
    .Y(_8047_)
);

OR2X2 _14283_ (
    .A(\datapath_1.ALUResult [14]),
    .B(_3671__bF$buf4),
    .Y(_3635_)
);

FILL FILL287280x64220 (
);

FILL FILL304760x113620 (
);

FILL FILL234840x118560 (
);

OR2X2 _15488_ (
    .A(_4440_),
    .B(_4441_),
    .Y(_4442_)
);

AND2X2 _15068_ (
    .A(_4048_),
    .B(_4055_),
    .Y(_4056_)
);

FILL FILL498560x167960 (
);

FILL FILL_0__16984_ (
);

FILL FILL_0__16564_ (
);

FILL FILL302480x187720 (
);

AND2X2 _8771_ (
    .A(_172_),
    .B(_171_),
    .Y(_135_[18])
);

FILL FILL251560x355680 (
);

FILL FILL21280x360620 (
);

FILL FILL_1__18776_ (
);

FILL FILL_1__13491_ (
);

OR2X2 _17634_ (
    .A(_6555_),
    .B(_6548_),
    .Y(_6556_)
);

FILL FILL_0__17349_ (
);

AND2X2 _17214_ (
    .A(_4160__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_6141_)
);

FILL FILL_0__12484_ (
);

FILL FILL201400x103740 (
);

FILL FILL_0__18710_ (
);

DFFSR _9976_ (
    .CLK(clk_bF$buf45),
    .D(_729_[4]),
    .Q(\datapath_1.regfile_1.regOut[12] [4]),
    .R(rst_bF$buf54),
    .S(vdd)
);

OR2X2 _9556_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .B(_596__bF$buf2),
    .Y(_576_)
);

OR2X2 _9136_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .B(_398__bF$buf0),
    .Y(_356_)
);

OR2X2 _18839_ (
    .A(_7709_),
    .B(_7742_),
    .Y(_7743_)
);

FILL FILL_0_BUFX2_insert560 (
);

AND2X2 _18419_ (
    .A(_6250__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_7329_)
);

FILL FILL_0_BUFX2_insert561 (
);

FILL FILL_0_BUFX2_insert562 (
);

FILL FILL_0_BUFX2_insert563 (
);

AND2X2 _13974_ (
    .A(_3344__bF$buf3),
    .B(gnd),
    .Y(_3397_)
);

FILL FILL_0__13689_ (
);

FILL FILL_0_BUFX2_insert564 (
);

AND2X2 _13554_ (
    .A(_3057_),
    .B(_3056_),
    .Y(_1_[21])
);

OR2X2 _13134_ (
    .A(_2157__bF$buf1),
    .B(_2685_),
    .Y(_2686_)
);

FILL FILL_0_BUFX2_insert566 (
);

FILL FILL_0_BUFX2_insert568 (
);

FILL FILL_0__14630_ (
);

FILL FILL_0__14210_ (
);

FILL FILL_1__9298_ (
);

FILL FILL8360x365560 (
);

FILL FILL505400x108680 (
);

OR2X2 _14759_ (
    .A(vdd),
    .B(_2_[1]),
    .Y(_3872_)
);

DFFSR _14339_ (
    .CLK(clk_bF$buf40),
    .D(_3606_[3]),
    .Q(ALUOut[3]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL145920x34580 (
);

FILL FILL158080x242060 (
);

FILL FILL_0__15835_ (
);

FILL FILL_0__15415_ (
);

AND2X2 _15700_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_4651_)
);

FILL FILL_0__10970_ (
);

FILL FILL_0__10550_ (
);

AND2X2 _18592_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_7499_)
);

AND2X2 _18172_ (
    .A(_6317__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_7086_)
);

FILL FILL_1__17627_ (
);

AND2X2 _10679_ (
    .A(_1144_),
    .B(_1143_),
    .Y(_1125_[9])
);

DFFSR _10259_ (
    .CLK(clk_bF$buf8),
    .D(_861_[29]),
    .Q(\datapath_1.regfile_1.regOut[14] [29]),
    .R(rst_bF$buf10),
    .S(vdd)
);

OR2X2 _16905_ (
    .A(_5836_),
    .B(_5829_),
    .Y(_5837_)
);

FILL FILL_0__11755_ (
);

OR2X2 _11620_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_1652__bF$buf3),
    .Y(_1632_)
);

FILL FILL_0__11335_ (
);

OR2X2 _11200_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_1454__bF$buf3),
    .Y(_1412_)
);

AND2X2 _19377_ (
    .A(_6216__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_8272_)
);

OR2X2 _14092_ (
    .A(_3498_),
    .B(_3495_),
    .Y(\datapath_1.alu_1.ALUInB [24])
);

FILL FILL367840x301340 (
);

DFFSR _8827_ (
    .CLK(clk_bF$buf5),
    .D(_135_[16]),
    .Q(\datapath_1.regfile_1.regOut[3] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

BUFX2 _8407_ (
    .A(_1_[15]),
    .Y(memoryAddress[15])
);

FILL FILL348840x138320 (
);

FILL FILL_1__13967_ (
);

FILL FILL503880x167960 (
);

AND2X2 _12825_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2390_)
);

OR2X2 _12405_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_2035_)
);

FILL FILL57000x271700 (
);

FILL FILL110200x128440 (
);

OR2X2 _15297_ (
    .A(_4253_),
    .B(_4250_),
    .Y(_4254_)
);

FILL FILL_0__13901_ (
);

FILL FILL_1__17380_ (
);

FILL FILL_1__8989_ (
);

FILL FILL209760x9880 (
);

DFFSR _8580_ (
    .CLK(clk_bF$buf59),
    .D(_3_[27]),
    .Q(\datapath_1.regfile_1.regOut[1] [27]),
    .R(rst_bF$buf25),
    .S(vdd)
);

FILL FILL270560x335920 (
);

FILL FILL105640x247000 (
);

FILL FILL180880x34580 (
);

FILL FILL196080x276640 (
);

FILL FILL_0__17998_ (
);

FILL FILL_0__17578_ (
);

OR2X2 _17863_ (
    .A(_6750_),
    .B(_6781_),
    .Y(_6782_)
);

AND2X2 _17443_ (
    .A(_6297__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_6368_)
);

AND2X2 _17023_ (
    .A(_4177__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_5953_)
);

FILL FILL369360x296400 (
);

FILL FILL501600x138320 (
);

AND2X2 _9785_ (
    .A(_688_),
    .B(_687_),
    .Y(_663_[12])
);

AND2X2 _9365_ (
    .A(_468_),
    .B(_467_),
    .Y(_465_[1])
);

FILL FILL_0__8620_ (
);

FILL FILL_0__10606_ (
);

OR2X2 _18648_ (
    .A(_7552_),
    .B(_7553_),
    .Y(_7554_)
);

AND2X2 _18228_ (
    .A(_6302__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_7141_)
);

AND2X2 _13783_ (
    .A(_3087__bF$buf0),
    .B(\datapath_1.ALUResult [27]),
    .Y(_3251_)
);

FILL FILL_0__13078_ (
);

XOR2X1 _13363_ (
    .A(_2189_),
    .B(_2901_),
    .Y(_2902_)
);

FILL FILL145160x247000 (
);

CLKBUF1 CLKBUF1_insert110 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf113)
);

CLKBUF1 CLKBUF1_insert111 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf112)
);

CLKBUF1 CLKBUF1_insert112 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf111)
);

FILL FILL104120x79040 (
);

CLKBUF1 CLKBUF1_insert113 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf110)
);

FILL FILL_0__9825_ (
);

CLKBUF1 CLKBUF1_insert114 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf109)
);

CLKBUF1 CLKBUF1_insert115 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf108)
);

CLKBUF1 CLKBUF1_insert116 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf107)
);

CLKBUF1 CLKBUF1_insert117 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf106)
);

CLKBUF1 CLKBUF1_insert118 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf105)
);

CLKBUF1 CLKBUF1_insert119 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf104)
);

FILL FILL366320x192660 (
);

DFFSR _14988_ (
    .CLK(clk_bF$buf12),
    .D(_3936_[7]),
    .Q(\datapath_1.mux_iord.din0 [7]),
    .R(rst_bF$buf91),
    .S(vdd)
);

OR2X2 _14568_ (
    .A(memoryOutData[23]),
    .B(_3803__bF$buf4),
    .Y(_3785_)
);

AND2X2 _14148_ (
    .A(_3543_),
    .B(_3542_),
    .Y(\datapath_1.mux_wd3.dout [1])
);

FILL FILL_1__16231_ (
);

FILL FILL335920x14820 (
);

FILL FILL_0__15224_ (
);

FILL FILL348840x365560 (
);

FILL FILL188480x291460 (
);

FILL FILL379240x59280 (
);

FILL FILL_1__17856_ (
);

DFFSR _10488_ (
    .CLK(clk_bF$buf69),
    .D(_993_[0]),
    .Q(\datapath_1.regfile_1.regOut[16] [0]),
    .R(rst_bF$buf76),
    .S(vdd)
);

OR2X2 _10068_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_837_)
);

FILL FILL_0__16849_ (
);

AND2X2 _16714_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_5649_)
);

FILL FILL_0__16429_ (
);

FILL FILL_0__11564_ (
);

AND2X2 _19186_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_8084_)
);

AND2X2 _8636_ (
    .A(_102_),
    .B(_101_),
    .Y(_69_[16])
);

FILL FILL252320x44460 (
);

FILL FILL_1__13356_ (
);

AND2X2 _17919_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_6837_)
);

OR2X2 _12634_ (
    .A(_2196_),
    .B(_2198_),
    .Y(_2199_)
);

FILL FILL_0__12349_ (
);

OR2X2 _12214_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .B(_1982__bF$buf1),
    .Y(_1928_)
);

FILL FILL427120x54340 (
);

FILL FILL_0__16182_ (
);

AND2X2 _13839_ (
    .A(_3292_),
    .B(_3291_),
    .Y(\datapath_1.alu_1.ALUInA [7])
);

NAND3X1 _13419_ (
    .A(_2383_),
    .B(_2500_),
    .C(_2389_),
    .Y(_2954_)
);

FILL FILL_1__15922_ (
);

FILL FILL_0__14915_ (
);

FILL FILL_0__17387_ (
);

AND2X2 _17672_ (
    .A(_6216__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_6593_)
);

AND2X2 _17252_ (
    .A(_4234__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_6179_)
);

FILL FILL91200x316160 (
);

DFFSR _9594_ (
    .CLK(clk_bF$buf102),
    .D(_531_[9]),
    .Q(\datapath_1.regfile_1.regOut[9] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

OR2X2 _9174_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_381_)
);

FILL FILL241680x370500 (
);

FILL FILL_0__10835_ (
);

FILL FILL_0__10415_ (
);

AND2X2 _10700_ (
    .A(_1158_),
    .B(_1157_),
    .Y(_1125_[16])
);

OR2X2 _18877_ (
    .A(_7779_),
    .B(_7776_),
    .Y(_7780_)
);

FILL FILL_0_BUFX2_insert940 (
);

FILL FILL_0_BUFX2_insert941 (
);

OR2X2 _18457_ (
    .A(_7362_),
    .B(_7365_),
    .Y(_7366_)
);

FILL FILL_0_BUFX2_insert942 (
);

AND2X2 _18037_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_6953_)
);

FILL FILL_0_BUFX2_insert943 (
);

FILL FILL_0_BUFX2_insert944 (
);

NOR2X1 _13592_ (
    .A(ALUOp[0]),
    .B(PCSource[1]),
    .Y(_3087_)
);

FILL FILL_0_BUFX2_insert946 (
);

AOI22X1 _13172_ (
    .A(_2720_),
    .B(_2379__bF$buf0),
    .C(_2593_),
    .D(_2721_),
    .Y(_2722_)
);

FILL FILL_0_BUFX2_insert948 (
);

FILL FILL_0__19113_ (
);

FILL FILL3040x261820 (
);

FILL FILL_0__9634_ (
);

OR2X2 _11905_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_1784__bF$buf4),
    .Y(_1782_)
);

AND2X2 _14797_ (
    .A(_3897_),
    .B(_3896_),
    .Y(_3870_[13])
);

FILL FILL385320x172900 (
);

AND2X2 _14377_ (
    .A(_3677_),
    .B(_3676_),
    .Y(_3672_[2])
);

FILL FILL_1__16880_ (
);

FILL FILL462080x54340 (
);

FILL FILL_0__15873_ (
);

FILL FILL_0__15453_ (
);

FILL FILL_0__15033_ (
);

FILL FILL408120x118560 (
);

FILL FILL252320x108680 (
);

FILL FILL47120x158080 (
);

OR2X2 _10297_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .B(_992__bF$buf0),
    .Y(_950_)
);

FILL FILL_1__17245_ (
);

OR2X2 _16943_ (
    .A(_5871_),
    .B(_5874_),
    .Y(_5875_)
);

AND2X2 _16523_ (
    .A(_4225__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_5461_)
);

OR2X2 _16103_ (
    .A(_5044_),
    .B(_5047_),
    .Y(_5048_)
);

OR2X2 _8865_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_215_)
);

BUFX2 _8445_ (
    .A(_2_[21]),
    .Y(memoryWriteData[21])
);

FILL FILL50920x192660 (
);

FILL FILL_1__13585_ (
);

AND2X2 _17728_ (
    .A(_6211__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_6649_)
);

OR2X2 _17308_ (
    .A(_6233_),
    .B(_6230_),
    .Y(_6234_)
);

OR2X2 _12863_ (
    .A(_2427_),
    .B(_2426_),
    .Y(_2428_)
);

FILL FILL_0__12578_ (
);

DFFSR _12443_ (
    .CLK(clk_bF$buf56),
    .D(_1983_[20]),
    .Q(\datapath_1.regfile_1.regOut[31] [20]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL_0__12158_ (
);

AND2X2 _12023_ (
    .A(_1840_),
    .B(_1839_),
    .Y(_1785_[27])
);

FILL FILL85120x79040 (
);

FILL FILL283480x306280 (
);

FILL FILL254600x197600 (
);

FILL FILL_0__8905_ (
);

FILL FILL237880x172900 (
);

AND2X2 _13648_ (
    .A(_3084__bF$buf1),
    .B(\datapath_1.PCJump [8]),
    .Y(_3135_)
);

XOR2X1 _13228_ (
    .A(_2214_),
    .B(_2774_),
    .Y(_2775_)
);

FILL FILL186960x340860 (
);

FILL FILL287280x227240 (
);

FILL FILL_0__14304_ (
);

FILL FILL497040x103740 (
);

OR2X2 _17481_ (
    .A(_6404_),
    .B(_6403_),
    .Y(_6405_)
);

FILL FILL_0__17196_ (
);

AND2X2 _17061_ (
    .A(_4130__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_5991_)
);

FILL FILL_0_CLKBUF1_insert170 (
);

FILL FILL_0_CLKBUF1_insert171 (
);

FILL FILL_0_CLKBUF1_insert172 (
);

FILL FILL_0__15929_ (
);

FILL FILL_0_CLKBUF1_insert174 (
);

FILL FILL_0_CLKBUF1_insert176 (
);

FILL FILL_0_CLKBUF1_insert178 (
);

FILL FILL_0__10224_ (
);

OR2X2 _18686_ (
    .A(_7590_),
    .B(_7591_),
    .Y(_7592_)
);

AND2X2 _18266_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_7178_)
);

FILL FILL_0__19342_ (
);

FILL FILL63080x88920 (
);

FILL FILL276640x74100 (
);

FILL FILL_0__11849_ (
);

FILL FILL_0__9023_ (
);

AND2X2 _11714_ (
    .A(_1674_),
    .B(_1673_),
    .Y(_1653_[10])
);

FILL FILL265240x281580 (
);

FILL FILL271320x222300 (
);

OR2X2 _14186_ (
    .A(\datapath_1.Data [14]),
    .B(_3605__bF$buf2),
    .Y(_3569_)
);

FILL FILL253080x74100 (
);

FILL FILL148960x123500 (
);

FILL FILL_0__15682_ (
);

AND2X2 _12919_ (
    .A(_2480_),
    .B(_2483_),
    .Y(_2484_)
);

FILL FILL_1_BUFX2_insert492 (
);

FILL FILL_1_BUFX2_insert494 (
);

FILL FILL_1_BUFX2_insert496 (
);

FILL FILL_1__17894_ (
);

FILL FILL438520x167960 (
);

FILL FILL66120x138320 (
);

AND2X2 _16752_ (
    .A(_4234__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_5687_)
);

FILL FILL_0__16467_ (
);

FILL FILL_0__16047_ (
);

OR2X2 _16332_ (
    .A(_5272_),
    .B(_5271_),
    .Y(_5273_)
);

FILL FILL234840x59280 (
);

OR2X2 _8674_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .B(_134__bF$buf3),
    .Y(_128_)
);

FILL FILL487160x192660 (
);

OR2X2 _17957_ (
    .A(_6873_),
    .B(_6870_),
    .Y(_6874_)
);

OR2X2 _17537_ (
    .A(_6445_),
    .B(_6460_),
    .Y(_6461_)
);

AND2X2 _17117_ (
    .A(_4234__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_6046_)
);

OR2X2 _12672_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2236_),
    .Y(_2237_)
);

FILL FILL_0__12387_ (
);

OR2X2 _12252_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_1953_)
);

FILL FILL_0__18613_ (
);

OR2X2 _9879_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_731_)
);

DFFSR _9459_ (
    .CLK(clk_bF$buf57),
    .D(_465_[3]),
    .Q(\datapath_1.regfile_1.regOut[8] [3]),
    .R(rst_bF$buf81),
    .S(vdd)
);

OR2X2 _9039_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_311_)
);

FILL FILL_0__8714_ (
);

OR2X2 _13877_ (
    .A(\datapath_1.a [20]),
    .B(_3342__bF$buf1),
    .Y(_3318_)
);

AND2X2 _13457_ (
    .A(_2989_),
    .B(_2918_),
    .Y(_2990_)
);

AND2X2 _13037_ (
    .A(_2591_),
    .B(_2594_),
    .Y(_2595_)
);

FILL FILL_0__14953_ (
);

FILL FILL_0__14533_ (
);

AND2X2 _17290_ (
    .A(_6215_),
    .B(_6201_),
    .Y(_6216_)
);

FILL FILL_0__9919_ (
);

FILL FILL349600x118560 (
);

FILL FILL_1__16745_ (
);

FILL FILL_1__16325_ (
);

FILL FILL_1__11880_ (
);

FILL FILL_1__11040_ (
);

FILL FILL_0__15318_ (
);

AND2X2 _15603_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_4556_)
);

FILL FILL_0__10033_ (
);

OR2X2 _18495_ (
    .A(_7403_),
    .B(_7400_),
    .Y(_7404_)
);

OR2X2 _18075_ (
    .A(_6986_),
    .B(_6989_),
    .Y(_6990_)
);

FILL FILL_0__19151_ (
);

FILL FILL453720x360620 (
);

FILL FILL197600x350740 (
);

FILL FILL16720x83980 (
);

FILL FILL_1__12245_ (
);

OR2X2 _16808_ (
    .A(_5741_),
    .B(_5734_),
    .Y(_5742_)
);

FILL FILL361000x74100 (
);

FILL FILL_0__9672_ (
);

OR2X2 _11943_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[28] [1]),
    .Y(_1787_)
);

FILL FILL294880x301340 (
);

DFFSR _11523_ (
    .CLK(clk_bF$buf57),
    .D(_1521_[3]),
    .Q(\datapath_1.regfile_1.regOut[24] [3]),
    .R(rst_bF$buf81),
    .S(vdd)
);

FILL FILL_0__11238_ (
);

OR2X2 _11103_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_1367_)
);

FILL FILL212040x301340 (
);

FILL FILL_0__15071_ (
);

NAND3X1 _12728_ (
    .A(_2282_),
    .B(\datapath_1.alu_1.ALUInA [16]),
    .C(_2292_),
    .Y(_2293_)
);

DFFSR _12308_ (
    .CLK(clk_bF$buf67),
    .D(_1917_[14]),
    .Q(\datapath_1.regfile_1.regOut[30] [14]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_0__16696_ (
);

AND2X2 _16981_ (
    .A(_4130__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_5912_)
);

AND2X2 _16561_ (
    .A(_4183__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_5499_)
);

FILL FILL_0__16276_ (
);

AND2X2 _16141_ (
    .A(_4167__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_5085_)
);

AND2X2 _8483_ (
    .A(_20_),
    .B(_19_),
    .Y(_3_[8])
);

FILL FILL_1__18068_ (
);

AND2X2 _17766_ (
    .A(_6282__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_6686_)
);

AND2X2 _17346_ (
    .A(_6220_),
    .B(_6201_),
    .Y(_6272_)
);

AND2X2 _12481_ (
    .A(_2058_),
    .B(_2072_),
    .Y(_2073_)
);

DFFSR _12061_ (
    .CLK(clk_bF$buf69),
    .D(_1785_[25]),
    .Q(\datapath_1.regfile_1.regOut[28] [25]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL30400x44460 (
);

FILL FILL345800x148200 (
);

FILL FILL_0__18842_ (
);

OR2X2 _9688_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .B(_662__bF$buf0),
    .Y(_644_)
);

OR2X2 _9268_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .B(_464__bF$buf1),
    .Y(_424_)
);

FILL FILL321480x54340 (
);

FILL FILL_1__11516_ (
);

FILL FILL_0__10929_ (
);

AND2X2 _13686_ (
    .A(_3089__bF$buf2),
    .B(gnd),
    .Y(_3168_)
);

NOR2X1 _13266_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2810_)
);

FILL FILL377720x123500 (
);

FILL FILL_0__19207_ (
);

FILL FILL_0__14762_ (
);

FILL FILL_0__9308_ (
);

FILL FILL_1__16974_ (
);

FILL FILL_0__15967_ (
);

OR2X2 _15832_ (
    .A(_4780_),
    .B(_4773_),
    .Y(_4781_)
);

FILL FILL_0__15547_ (
);

AND2X2 _15412_ (
    .A(_4183__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_4368_)
);

FILL FILL_0__10262_ (
);

FILL FILL202920x350740 (
);

FILL FILL_0__19380_ (
);

FILL FILL94240x370500 (
);

FILL FILL385320x335920 (
);

FILL FILL129960x306280 (
);

FILL FILL320720x247000 (
);

AND2X2 _16617_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_5554_)
);

FILL FILL326040x321100 (
);

FILL FILL_0__11887_ (
);

OR2X2 _11752_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .B(_1718__bF$buf3),
    .Y(_1700_)
);

FILL FILL_0__11467_ (
);

FILL FILL_0__9061_ (
);

FILL FILL_0__11047_ (
);

OR2X2 _11332_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .B(_1520__bF$buf3),
    .Y(_1480_)
);

AND2X2 _19089_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_7989_)
);

DFFSR _8959_ (
    .CLK(clk_bF$buf19),
    .D(_201_[19]),
    .Q(\datapath_1.regfile_1.regOut[4] [19]),
    .R(rst_bF$buf13),
    .S(vdd)
);

OR2X2 _8539_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .B(_68__bF$buf3),
    .Y(_58_)
);

FILL FILL256120x326040 (
);

FILL FILL197600x59280 (
);

OR2X2 _9900_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_745_)
);

NOR2X1 _12957_ (
    .A(_2519_),
    .B(_2517_),
    .Y(_2520_)
);

FILL FILL_1_BUFX2_insert872 (
);

OR2X2 _12537_ (
    .A(_2126_),
    .B(_2124_),
    .Y(_2127_)
);

FILL FILL_1_BUFX2_insert874 (
);

OR2X2 _12117_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_1883_)
);

FILL FILL_1_BUFX2_insert876 (
);

FILL FILL4560x143260 (
);

FILL FILL_0__13613_ (
);

FILL FILL209000x64220 (
);

OR2X2 _16790_ (
    .A(_5723_),
    .B(_5722_),
    .Y(_5724_)
);

OR2X2 _16370_ (
    .A(_5310_),
    .B(_5309_),
    .Y(_5311_)
);

FILL FILL424080x167960 (
);

FILL FILL199880x54340 (
);

FILL FILL_1__18297_ (
);

BUFX2 BUFX2_insert540 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf99)
);

BUFX2 BUFX2_insert541 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf98)
);

BUFX2 BUFX2_insert542 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf97)
);

BUFX2 BUFX2_insert543 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf96)
);

AND2X2 _17995_ (
    .A(_6911_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd1 [9])
);

BUFX2 BUFX2_insert544 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf95)
);

BUFX2 BUFX2_insert545 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf94)
);

AND2X2 _17575_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_6498_)
);

FILL FILL152760x24700 (
);

AND2X2 _17155_ (
    .A(_4154__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_6083_)
);

BUFX2 BUFX2_insert546 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf93)
);

BUFX2 BUFX2_insert547 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf92)
);

BUFX2 BUFX2_insert548 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf91)
);

BUFX2 BUFX2_insert549 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf90)
);

AND2X2 _12290_ (
    .A(_1978_),
    .B(_1977_),
    .Y(_1917_[30])
);

FILL FILL_0__18231_ (
);

FILL FILL437000x14820 (
);

AND2X2 _9497_ (
    .A(_536_),
    .B(_535_),
    .Y(_531_[2])
);

DFFSR _9077_ (
    .CLK(clk_bF$buf37),
    .D(_267_[8]),
    .Q(\datapath_1.regfile_1.regOut[5] [8]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_1__11325_ (
);

FILL FILL_0__8752_ (
);

FILL FILL_0__10738_ (
);

FILL FILL_0__10318_ (
);

OR2X2 _10603_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_1124__bF$buf4),
    .Y(_1114_)
);

FILL FILL_0_BUFX2_insert60 (
);

FILL FILL_0_BUFX2_insert61 (
);

FILL FILL_0_BUFX2_insert62 (
);

FILL FILL_0_BUFX2_insert64 (
);

FILL FILL_0_BUFX2_insert66 (
);

OR2X2 _13495_ (
    .A(IorD_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [2]),
    .Y(_3018_)
);

XOR2X1 _13075_ (
    .A(_2613_),
    .B(_2617_),
    .Y(_2631_)
);

FILL FILL_0_BUFX2_insert68 (
);

FILL FILL_0__19436_ (
);

FILL FILL_0__19016_ (
);

AND2X2 _19301_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_8197_)
);

FILL FILL_0__14571_ (
);

FILL FILL504640x217360 (
);

FILL FILL_0__9957_ (
);

DFFSR _11808_ (
    .CLK(clk_bF$buf32),
    .D(_1653_[30]),
    .Q(\datapath_1.regfile_1.regOut[26] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL_0__9117_ (
);

FILL FILL405080x113620 (
);

FILL FILL156560x24700 (
);

FILL FILL383800x39520 (
);

FILL FILL_1__16363_ (
);

FILL FILL29640x281580 (
);

OR2X2 _15641_ (
    .A(_4577_),
    .B(_4592_),
    .Y(_4593_)
);

OR2X2 _15221_ (
    .A(_4176_),
    .B(_4178_),
    .Y(_4179_)
);

FILL FILL12160x365560 (
);

FILL FILL205960x34580 (
);

FILL FILL333640x286520 (
);

AND2X2 _16846_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_5779_)
);

AND2X2 _16426_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_5366_)
);

AND2X2 _16006_ (
    .A(_4197__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_4952_)
);

AND2X2 _11981_ (
    .A(_1812_),
    .B(_1811_),
    .Y(_1785_[13])
);

FILL FILL_0__11696_ (
);

FILL FILL_0__9290_ (
);

AND2X2 _11561_ (
    .A(_1592_),
    .B(_1591_),
    .Y(_1587_[2])
);

DFFSR _11141_ (
    .CLK(clk_bF$buf21),
    .D(_1323_[8]),
    .Q(\datapath_1.regfile_1.regOut[21] [8]),
    .R(rst_bF$buf4),
    .S(vdd)
);

FILL FILL_0__17502_ (
);

FILL FILL269040x365560 (
);

AND2X2 _8768_ (
    .A(_170_),
    .B(_169_),
    .Y(_135_[17])
);

FILL FILL356440x370500 (
);

FILL FILL384560x103740 (
);

NAND2X1 _12766_ (
    .A(\datapath_1.alu_1.ALUInA [24]),
    .B(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2331_)
);

OR2X2 _12346_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .B(_2048__bF$buf4),
    .Y(_1996_)
);

FILL FILL_0__18707_ (
);

FILL FILL_0__13842_ (
);

FILL FILL_0__13422_ (
);

FILL FILL491720x54340 (
);

FILL FILL300200x271700 (
);

FILL FILL_1__15214_ (
);

FILL FILL299440x187720 (
);

OR2X2 _14912_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [9]),
    .Y(_3954_)
);

FILL FILL_0__14207_ (
);

FILL FILL437000x103740 (
);

OR2X2 _17384_ (
    .A(_6201_),
    .B(_6309_),
    .Y(_6310_)
);

FILL FILL_0__18880_ (
);

FILL FILL_0__18460_ (
);

FILL FILL_1__16839_ (
);

FILL FILL_0__8981_ (
);

FILL FILL_0__10547_ (
);

AND2X2 _10832_ (
    .A(_1226_),
    .B(_1225_),
    .Y(_1191_[17])
);

AND2X2 _10412_ (
    .A(_1006_),
    .B(_1005_),
    .Y(_993_[6])
);

AND2X2 _18589_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_7496_)
);

OR2X2 _18169_ (
    .A(_7079_),
    .B(_7082_),
    .Y(_7083_)
);

DFFSR _19530_ (
    .CLK(clk_bF$buf18),
    .D(_8320_[7]),
    .Q(\datapath_1.regfile_1.regOut[0] [7]),
    .R(rst_bF$buf107),
    .S(vdd)
);

OR2X2 _19110_ (
    .A(_8007_),
    .B(_8008_),
    .Y(_8009_)
);

FILL FILL_0__14380_ (
);

FILL FILL_0__9766_ (
);

FILL FILL348840x251940 (
);

OR2X2 _11617_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .B(_1652__bF$buf0),
    .Y(_1630_)
);

FILL FILL449160x138320 (
);

AND2X2 _14089_ (
    .A(_3350__bF$buf1),
    .B(_2_[24]),
    .Y(_3496_)
);

FILL FILL248520x345800 (
);

FILL FILL278920x256880 (
);

AND2X2 _15870_ (
    .A(_4181__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_4818_)
);

FILL FILL_0__15585_ (
);

FILL FILL_0__15165_ (
);

AND2X2 _15450_ (
    .A(_4160__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_4405_)
);

INVX1 _15030_ (
    .A(\datapath_1.a3 [2]),
    .Y(_4019_)
);

FILL FILL475000x271700 (
);

FILL FILL466640x148200 (
);

FILL FILL106400x34580 (
);

FILL FILL297160x370500 (
);

OR2X2 _16655_ (
    .A(_5589_),
    .B(_5590_),
    .Y(_5591_)
);

OR2X2 _16235_ (
    .A(_5176_),
    .B(_5177_),
    .Y(_5178_)
);

FILL FILL38760x69160 (
);

FILL FILL105640x360620 (
);

DFFSR _11790_ (
    .CLK(clk_bF$buf103),
    .D(_1653_[12]),
    .Q(\datapath_1.regfile_1.regOut[26] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

OR2X2 _11370_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_1505_)
);

FILL FILL_0__11085_ (
);

FILL FILL_0__17731_ (
);

FILL FILL_0__17311_ (
);

OR2X2 _8997_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_283_)
);

DFFSR _8577_ (
    .CLK(clk_bF$buf35),
    .D(_3_[24]),
    .Q(\datapath_1.regfile_1.regOut[1] [24]),
    .R(rst_bF$buf6),
    .S(vdd)
);

FILL FILL288040x345800 (
);

FILL FILL_1__10825_ (
);

AND2X2 _12995_ (
    .A(_2555_),
    .B(_2553_),
    .Y(_2556_)
);

OR2X2 _12575_ (
    .A(vdd),
    .B(\control_1.reg_state.dout [1]),
    .Y(_2147_)
);

AND2X2 _12155_ (
    .A(_1908_),
    .B(_1907_),
    .Y(_1851_[28])
);

AND2X2 _18801_ (
    .A(_6293__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_7705_)
);

FILL FILL259920x202540 (
);

FILL FILL312360x44460 (
);

FILL FILL244720x19760 (
);

FILL FILL_0__8617_ (
);

FILL FILL_1__9680_ (
);

BUFX2 BUFX2_insert1100 (
    .A(_1322_),
    .Y(_1322__bF$buf4)
);

FILL FILL253840x355680 (
);

BUFX2 BUFX2_insert1101 (
    .A(_1322_),
    .Y(_1322__bF$buf3)
);

BUFX2 BUFX2_insert1102 (
    .A(_1322_),
    .Y(_1322__bF$buf2)
);

BUFX2 BUFX2_insert1103 (
    .A(_1322_),
    .Y(_1322__bF$buf1)
);

FILL FILL23560x360620 (
);

BUFX2 BUFX2_insert1104 (
    .A(_1322_),
    .Y(_1322__bF$buf0)
);

BUFX2 BUFX2_insert1105 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf4 )
);

BUFX2 BUFX2_insert1106 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf3 )
);

BUFX2 BUFX2_insert1107 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf2 )
);

FILL FILL_1__15863_ (
);

FILL FILL_1__15443_ (
);

BUFX2 BUFX2_insert1108 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf1 )
);

BUFX2 BUFX2_insert1109 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf0 )
);

OR2X2 _14721_ (
    .A(\datapath_1.rd1 [31]),
    .B(_3869__bF$buf2),
    .Y(_3867_)
);

FILL FILL_0__14436_ (
);

FILL FILL_0__14016_ (
);

OR2X2 _14301_ (
    .A(\datapath_1.ALUResult [20]),
    .B(_3671__bF$buf0),
    .Y(_3647_)
);

BUFX2 BUFX2_insert920 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf2 )
);

BUFX2 BUFX2_insert921 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf1 )
);

BUFX2 BUFX2_insert922 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf0 )
);

BUFX2 BUFX2_insert923 (
    .A(_3342_),
    .Y(_3342__bF$buf4)
);

BUFX2 BUFX2_insert924 (
    .A(_3342_),
    .Y(_3342__bF$buf3)
);

BUFX2 BUFX2_insert925 (
    .A(_3342_),
    .Y(_3342__bF$buf2)
);

BUFX2 BUFX2_insert926 (
    .A(_3342_),
    .Y(_3342__bF$buf1)
);

AND2X2 _17193_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_6121_)
);

BUFX2 BUFX2_insert927 (
    .A(_3342_),
    .Y(_3342__bF$buf0)
);

BUFX2 BUFX2_insert928 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf4 )
);

BUFX2 BUFX2_insert929 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf3 )
);

OR2X2 _15926_ (
    .A(_4870_),
    .B(_4873_),
    .Y(_4874_)
);

AND2X2 _15506_ (
    .A(_4241__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_4460_)
);

FILL FILL_0__8790_ (
);

FILL FILL_0__10356_ (
);

DFFSR _10641_ (
    .CLK(clk_bF$buf35),
    .D(_1059_[24]),
    .Q(\datapath_1.regfile_1.regOut[17] [24]),
    .R(rst_bF$buf67),
    .S(vdd)
);

OR2X2 _10221_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_919_)
);

OR2X2 _18398_ (
    .A(_7306_),
    .B(_7307_),
    .Y(_7308_)
);

FILL FILL316160x44460 (
);

FILL FILL_0__19474_ (
);

FILL FILL_0__19054_ (
);

FILL FILL231800x4940 (
);

FILL FILL_1__12568_ (
);

AND2X2 _11846_ (
    .A(_1742_),
    .B(_1741_),
    .Y(_1719_[11])
);

AND2X2 _11426_ (
    .A(_1522_),
    .B(_1585_),
    .Y(_1521_[0])
);

DFFSR _11006_ (
    .CLK(clk_bF$buf111),
    .D(_1257_[2]),
    .Q(\datapath_1.regfile_1.regOut[20] [2]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL498560x350740 (
);

FILL FILL321480x212420 (
);

FILL FILL_0__15394_ (
);

FILL FILL361000x321100 (
);

FILL FILL_1__14714_ (
);

FILL FILL177080x158080 (
);

FILL FILL_0__13707_ (
);

FILL FILL_1__17186_ (
);

AND2X2 _16884_ (
    .A(_4135__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [25]),
    .Y(_5817_)
);

OR2X2 _16464_ (
    .A(_5402_),
    .B(_5399_),
    .Y(_5403_)
);

AND2X2 _16044_ (
    .A(_4203__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_4990_)
);

FILL FILL_0__17960_ (
);

FILL FILL_1__10214_ (
);

FILL FILL374680x44460 (
);

FILL FILL236360x296400 (
);

OR2X2 _17669_ (
    .A(_6557_),
    .B(_6590_),
    .Y(_6591_)
);

AND2X2 _17249_ (
    .A(_4200__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_6176_)
);

FILL FILL126920x64220 (
);

OR2X2 _12384_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_2021_)
);

FILL FILL_0__12099_ (
);

FILL FILL395200x340860 (
);

FILL FILL_0__18745_ (
);

FILL FILL283480x19760 (
);

FILL FILL_0__18325_ (
);

OR2X2 _18610_ (
    .A(_7502_),
    .B(_7516_),
    .Y(_7517_)
);

FILL FILL_0__13460_ (
);

FILL FILL_0__13040_ (
);

FILL FILL120080x14820 (
);

FILL FILL_0__8426_ (
);

FILL FILL298680x182780 (
);

FILL FILL234080x83980 (
);

AND2X2 _13589_ (
    .A(_3083_),
    .B(PCSource[1]),
    .Y(_3084_)
);

FILL FILL123120x79040 (
);

AOI22X1 _13169_ (
    .A(_2718_),
    .B(_2504_),
    .C(_2548_),
    .D(_2717_),
    .Y(_2719_)
);

FILL FILL107920x247000 (
);

FILL FILL_0__14665_ (
);

AND2X2 _14950_ (
    .A(_3979_),
    .B(_3978_),
    .Y(_3936_[21])
);

AND2X2 _14530_ (
    .A(_3759_),
    .B(_3758_),
    .Y(_3738_[10])
);

AND2X2 _14110_ (
    .A(_3350__bF$buf1),
    .B(_2_[27]),
    .Y(_3514_)
);

OR2X2 _15735_ (
    .A(_4678_),
    .B(_4685_),
    .Y(_4686_)
);

OR2X2 _15315_ (
    .A(_4270_),
    .B(_4271_),
    .Y(_4272_)
);

FILL FILL_0__10585_ (
);

OR2X2 _10870_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .B(_1256__bF$buf0),
    .Y(_1252_)
);

OR2X2 _10450_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .B(_1058__bF$buf2),
    .Y(_1032_)
);

FILL FILL_0__10165_ (
);

OR2X2 _10030_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .B(_860__bF$buf0),
    .Y(_812_)
);

BUFX2 BUFX2_insert70 (
    .A(_4214_),
    .Y(_4214__bF$buf4)
);

BUFX2 BUFX2_insert71 (
    .A(_4214_),
    .Y(_4214__bF$buf3)
);

BUFX2 BUFX2_insert72 (
    .A(_4214_),
    .Y(_4214__bF$buf2)
);

BUFX2 BUFX2_insert73 (
    .A(_4214_),
    .Y(_4214__bF$buf1)
);

BUFX2 BUFX2_insert74 (
    .A(_4214_),
    .Y(_4214__bF$buf0)
);

FILL FILL_0__16811_ (
);

BUFX2 BUFX2_insert75 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf4 )
);

BUFX2 BUFX2_insert76 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf3 )
);

BUFX2 BUFX2_insert77 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf2 )
);

BUFX2 BUFX2_insert78 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf1 )
);

FILL FILL224960x256880 (
);

BUFX2 BUFX2_insert79 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf0 )
);

FILL FILL_0__19283_ (
);

FILL FILL34200x370500 (
);

FILL FILL_1__12377_ (
);

FILL FILL503880x350740 (
);

FILL FILL368600x192660 (
);

FILL FILL_1__18603_ (
);

DFFSR _11655_ (
    .CLK(clk_bF$buf14),
    .D(_1587_[6]),
    .Q(\datapath_1.regfile_1.regOut[25] [6]),
    .R(rst_bF$buf8),
    .S(vdd)
);

OR2X2 _11235_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_1435_)
);

FILL FILL124640x88920 (
);

FILL FILL110200x311220 (
);

FILL FILL_0__12731_ (
);

AND2X2 _9803_ (
    .A(_700_),
    .B(_699_),
    .Y(_663_[18])
);

FILL FILL336680x74100 (
);

FILL FILL22040x64220 (
);

FILL FILL_1__14523_ (
);

FILL FILL_1__14103_ (
);

FILL FILL_0__13936_ (
);

FILL FILL388360x321100 (
);

AND2X2 _13801_ (
    .A(_3081__bF$buf1),
    .B(ALUOut[30]),
    .Y(_3266_)
);

OR2X2 _16693_ (
    .A(_5627_),
    .B(_5628_),
    .Y(_5629_)
);

AND2X2 _16273_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_5215_)
);

FILL FILL_1__15728_ (
);

FILL FILL_1__15308_ (
);

FILL FILL_1__10023_ (
);

FILL FILL326040x281580 (
);

AND2X2 _17898_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_6816_)
);

OR2X2 _17478_ (
    .A(_6401_),
    .B(_6400_),
    .Y(_6402_)
);

AND2X2 _17058_ (
    .A(_4200__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_5988_)
);

DFFSR _12193_ (
    .CLK(clk_bF$buf91),
    .D(_1851_[28]),
    .Q(\datapath_1.regfile_1.regOut[29] [28]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL_0__18974_ (
);

FILL FILL_0__18554_ (
);

FILL FILL_0__18134_ (
);

FILL FILL262200x227240 (
);

FILL FILL_1__11228_ (
);

FILL FILL_0__8655_ (
);

OR2X2 _10926_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_1269_)
);

DFFSR _10506_ (
    .CLK(clk_bF$buf84),
    .D(_993_[18]),
    .Q(\datapath_1.regfile_1.regOut[16] [18]),
    .R(rst_bF$buf47),
    .S(vdd)
);

AND2X2 _13398_ (
    .A(_2934_),
    .B(_2922_),
    .Y(_2935_)
);

FILL FILL_1__15481_ (
);

AND2X2 _19204_ (
    .A(_6326__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_8102_)
);

FILL FILL_0__14894_ (
);

FILL FILL_0__14054_ (
);

FILL FILL427880x113620 (
);

FILL FILL207480x197600 (
);

FILL FILL396720x79040 (
);

FILL FILL412680x375440 (
);

OR2X2 _15964_ (
    .A(_4909_),
    .B(_4910_),
    .Y(_4911_)
);

FILL FILL_0__15679_ (
);

OR2X2 _15544_ (
    .A(_4497_),
    .B(_4482_),
    .Y(_4498_)
);

FILL FILL_0__15259_ (
);

AND2X2 _15124_ (
    .A(_4029_),
    .B(_4101_),
    .Y(\datapath_1.regfile_1.regEn [12])
);

FILL FILL_0__10394_ (
);

FILL FILL66120x251940 (
);

FILL FILL_0__16200_ (
);

FILL FILL5320x261820 (
);

AND2X2 _16749_ (
    .A(_4130__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_5684_)
);

OR2X2 _16329_ (
    .A(_5269_),
    .B(_5262_),
    .Y(_5270_)
);

FILL FILL387600x172900 (
);

OR2X2 _11884_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .B(_1784__bF$buf2),
    .Y(_1768_)
);

FILL FILL_0__11599_ (
);

FILL FILL_0__9193_ (
);

OR2X2 _11464_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_1586__bF$buf0),
    .Y(_1548_)
);

FILL FILL_0__11179_ (
);

OR2X2 _11044_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .B(_1388__bF$buf2),
    .Y(_1328_)
);

FILL FILL_0__17825_ (
);

FILL FILL_0__12960_ (
);

FILL FILL_0__12540_ (
);

FILL FILL_0__12120_ (
);

FILL FILL341240x153140 (
);

FILL FILL_1__10919_ (
);

FILL FILL378480x276640 (
);

DFFSR _9612_ (
    .CLK(clk_bF$buf66),
    .D(_531_[27]),
    .Q(\datapath_1.regfile_1.regOut[9] [27]),
    .R(rst_bF$buf80),
    .S(vdd)
);

OR2X2 _12669_ (
    .A(_2233_),
    .B(_2223_),
    .Y(_2234_)
);

OR2X2 _12249_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_1951_)
);

FILL FILL_1__14332_ (
);

FILL FILL395960x286520 (
);

FILL FILL472720x232180 (
);

FILL FILL_0__13325_ (
);

OR2X2 _13610_ (
    .A(_3102_),
    .B(_3101_),
    .Y(_3103_)
);

AND2X2 _16082_ (
    .A(_4230__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_5027_)
);

FILL FILL_1__15957_ (
);

FILL FILL32680x227240 (
);

AND2X2 _14815_ (
    .A(_3909_),
    .B(_3908_),
    .Y(_3870_[19])
);

FILL FILL505400x335920 (
);

OR2X2 _17287_ (
    .A(_6207_),
    .B(_6212_),
    .Y(_6213_)
);

FILL FILL285760x306280 (
);

FILL FILL427880x340860 (
);

FILL FILL_0__18783_ (
);

FILL FILL_0__8884_ (
);

FILL FILL_0__8464_ (
);

OR2X2 _10735_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .B(_1190__bF$buf0),
    .Y(_1182_)
);

OR2X2 _10315_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .B(_992__bF$buf3),
    .Y(_962_)
);

FILL FILL220400x316160 (
);

FILL FILL_0__11811_ (
);

FILL FILL499320x103740 (
);

OR2X2 _19433_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_8324_)
);

FILL FILL_0__19148_ (
);

OR2X2 _19013_ (
    .A(_7913_),
    .B(_7912_),
    .Y(_7914_)
);

FILL FILL158080x335920 (
);

FILL FILL_0__14283_ (
);

FILL FILL272080x74100 (
);

FILL FILL408120x301340 (
);

FILL FILL_0__9249_ (
);

FILL FILL175560x345800 (
);

AND2X2 _15773_ (
    .A(_4200__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_4723_)
);

FILL FILL_0__15488_ (
);

OR2X2 _15353_ (
    .A(_4309_),
    .B(_4278_),
    .Y(_4310_)
);

FILL FILL408880x54340 (
);

FILL FILL267520x281580 (
);

AND2X2 _16978_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_5909_)
);

OR2X2 _16558_ (
    .A(_5495_),
    .B(_5494_),
    .Y(_5496_)
);

AND2X2 _16138_ (
    .A(_4175__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_5082_)
);

FILL FILL273600x222300 (
);

AND2X2 _11693_ (
    .A(_1660_),
    .B(_1659_),
    .Y(_1653_[3])
);

DFFSR _11273_ (
    .CLK(clk_bF$buf95),
    .D(_1389_[11]),
    .Q(\datapath_1.regfile_1.regOut[22] [11]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL21280x29640 (
);

FILL FILL127680x266760 (
);

FILL FILL_0__17214_ (
);

FILL FILL9120x301340 (
);

OR2X2 _9841_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .B(_728__bF$buf4),
    .Y(_726_)
);

OR2X2 _9421_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .B(_530__bF$buf3),
    .Y(_506_)
);

OR2X2 _9001_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .B(_332__bF$buf3),
    .Y(_286_)
);

AND2X2 _12898_ (
    .A(_2462_),
    .B(_2278_),
    .Y(_2463_)
);

OAI21X1 _12478_ (
    .A(_2070_),
    .B(_2068_),
    .C(_2055_),
    .Y(_2071_)
);

DFFSR _12058_ (
    .CLK(clk_bF$buf74),
    .D(_1785_[22]),
    .Q(\datapath_1.regfile_1.regOut[28] [22]),
    .R(rst_bF$buf47),
    .S(vdd)
);

FILL FILL_0__18839_ (
);

OR2X2 _18704_ (
    .A(_7609_),
    .B(_7608_),
    .Y(_7610_)
);

FILL FILL_0__18419_ (
);

FILL FILL_0__13974_ (
);

FILL FILL_0__13554_ (
);

FILL FILL_0__13134_ (
);

FILL FILL_1__9583_ (
);

FILL FILL446120x335920 (
);

DFFSR _14624_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[30]),
    .Q(\control_1.op [4]),
    .R(rst_bF$buf100),
    .S(vdd)
);

OR2X2 _14204_ (
    .A(\datapath_1.Data [20]),
    .B(_3605__bF$buf4),
    .Y(_3581_)
);

OR2X2 _17096_ (
    .A(_6021_),
    .B(_6024_),
    .Y(_6025_)
);

FILL FILL389120x286520 (
);

FILL FILL_0__15700_ (
);

FILL FILL_0__18172_ (
);

FILL FILL161120x316160 (
);

FILL FILL303240x350740 (
);

FILL FILL_1__11686_ (
);

AND2X2 _15829_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_4778_)
);

FILL FILL504640x103740 (
);

AND2X2 _15409_ (
    .A(_4200__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_4365_)
);

FILL FILL85880x360620 (
);

AND2X2 _10964_ (
    .A(_1294_),
    .B(_1293_),
    .Y(_1257_[18])
);

FILL FILL_0__10679_ (
);

AND2X2 _10544_ (
    .A(_1074_),
    .B(_1073_),
    .Y(_1059_[7])
);

DFFSR _10124_ (
    .CLK(clk_bF$buf101),
    .D(_795_[23]),
    .Q(\datapath_1.regfile_1.regOut[13] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL66880x197600 (
);

FILL FILL_0__11620_ (
);

FILL FILL_0__11200_ (
);

AND2X2 _19242_ (
    .A(_6221__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_8139_)
);

FILL FILL151240x261820 (
);

FILL FILL_0__9058_ (
);

OR2X2 _11749_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_1718__bF$buf3),
    .Y(_1698_)
);

OR2X2 _11329_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .B(_1520__bF$buf4),
    .Y(_1478_)
);

FILL FILL_1__13832_ (
);

FILL FILL_0__12825_ (
);

FILL FILL_0__12405_ (
);

FILL FILL333640x172900 (
);

AND2X2 _15582_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_4535_)
);

NAND3X1 _15162_ (
    .A(_4030_),
    .B(\datapath_1.a3 [4]),
    .C(_4031_),
    .Y(_4124_)
);

FILL FILL282720x340860 (
);

FILL FILL_1__8434_ (
);

OR2X2 _16787_ (
    .A(_5719_),
    .B(_5720_),
    .Y(_5721_)
);

OR2X2 _16367_ (
    .A(_5304_),
    .B(_5307_),
    .Y(_5308_)
);

FILL FILL214320x301340 (
);

OR2X2 _11082_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_1353_)
);

FILL FILL_1__9639_ (
);

FILL FILL_0__17863_ (
);

FILL FILL_0__17443_ (
);

FILL FILL_0__17023_ (
);

FILL FILL240160x242060 (
);

FILL FILL_1__10957_ (
);

AND2X2 _9650_ (
    .A(_618_),
    .B(_617_),
    .Y(_597_[10])
);

OR2X2 _9230_ (
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .Y(_463_)
);

FILL FILL272840x29640 (
);

FILL FILL310080x103740 (
);

AND2X2 _12287_ (
    .A(_1976_),
    .B(_1975_),
    .Y(_1917_[29])
);

FILL FILL_0__18648_ (
);

OR2X2 _18933_ (
    .A(_7827_),
    .B(_7834_),
    .Y(_7835_)
);

OR2X2 _18513_ (
    .A(_7390_),
    .B(_7421_),
    .Y(_7422_)
);

FILL FILL_0__13783_ (
);

FILL FILL240160x108680 (
);

FILL FILL_0__8749_ (
);

FILL FILL26600x227240 (
);

DFFSR _14853_ (
    .CLK(clk_bF$buf94),
    .D(_3870_[1]),
    .Q(_2_[1]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL174800x128440 (
);

FILL FILL_0__14148_ (
);

OR2X2 _14433_ (
    .A(memoryOutData[21]),
    .B(_3737__bF$buf2),
    .Y(_3715_)
);

AND2X2 _14013_ (
    .A(_3352__bF$buf1),
    .B(\datapath_1.PCJump [13]),
    .Y(_3431_)
);

FILL FILL280440x202540 (
);

FILL FILL155800x286520 (
);

FILL FILL430160x365560 (
);

FILL FILL434720x93860 (
);

FILL FILL_1__11075_ (
);

OR2X2 _15638_ (
    .A(_4589_),
    .B(_4588_),
    .Y(_4590_)
);

AND2X2 _15218_ (
    .A(_4175__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_4176_)
);

FILL FILL_1__17721_ (
);

DFFSR _10773_ (
    .CLK(clk_bF$buf66),
    .D(_1125_[27]),
    .Q(\datapath_1.regfile_1.regOut[18] [27]),
    .R(rst_bF$buf69),
    .S(vdd)
);

FILL FILL_0__10068_ (
);

OR2X2 _10353_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_987_)
);

FILL FILL_0__16714_ (
);

AND2X2 _19471_ (
    .A(_8349_),
    .B(_8348_),
    .Y(_8320_[14])
);

FILL FILL_0__19186_ (
);

OR2X2 _19051_ (
    .A(_7942_),
    .B(_7950_),
    .Y(_7951_)
);

AND2X2 _8921_ (
    .A(_252_),
    .B(_251_),
    .Y(_201_[25])
);

AND2X2 _8501_ (
    .A(_32_),
    .B(_31_),
    .Y(_3_[14])
);

AND2X2 _11978_ (
    .A(_1810_),
    .B(_1809_),
    .Y(_1785_[12])
);

AND2X2 _11558_ (
    .A(_1590_),
    .B(_1589_),
    .Y(_1587_[1])
);

DFFSR _11138_ (
    .CLK(clk_bF$buf68),
    .D(_1323_[5]),
    .Q(\datapath_1.regfile_1.regOut[21] [5]),
    .R(rst_bF$buf40),
    .S(vdd)
);

FILL FILL_1__13221_ (
);

FILL FILL_0__17919_ (
);

FILL FILL_0__12214_ (
);

OR2X2 _15391_ (
    .A(_4345_),
    .B(_4346_),
    .Y(_4347_)
);

FILL FILL9880x247000 (
);

OR2X2 _9706_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .B(_662__bF$buf4),
    .Y(_656_)
);

FILL FILL204440x256880 (
);

FILL FILL_0__13839_ (
);

FILL FILL_0__13419_ (
);

AND2X2 _13704_ (
    .A(_3084__bF$buf3),
    .B(\datapath_1.PCJump [16]),
    .Y(_3183_)
);

AND2X2 _16596_ (
    .A(_4172__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_5533_)
);

AND2X2 _16176_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_5120_)
);

FILL FILL_1__9028_ (
);

FILL FILL_0__17672_ (
);

FILL FILL_0__17252_ (
);

FILL FILL_1__10346_ (
);

OR2X2 _14909_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [8]),
    .Y(_3952_)
);

FILL FILL131480x74100 (
);

FILL FILL_1__19464_ (
);

OR2X2 _12096_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_1869_)
);

FILL FILL_1__19044_ (
);

AND2X2 _18742_ (
    .A(_6238__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_7647_)
);

AND2X2 _18322_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_7233_)
);

FILL FILL_0__18037_ (
);

FILL FILL_0__13592_ (
);

FILL FILL_0__13172_ (
);

AND2X2 _10829_ (
    .A(_1224_),
    .B(_1223_),
    .Y(_1191_[16])
);

FILL FILL124640x232180 (
);

AND2X2 _10409_ (
    .A(_1004_),
    .B(_1003_),
    .Y(_993_[5])
);

FILL FILL33440x0 (
);

DFFSR _19527_ (
    .CLK(clk_bF$buf73),
    .D(_8320_[4]),
    .Q(\datapath_1.regfile_1.regOut[0] [4]),
    .R(rst_bF$buf39),
    .S(vdd)
);

OR2X2 _19107_ (
    .A(_8002_),
    .B(_8005_),
    .Y(_8006_)
);

FILL FILL_0__14797_ (
);

AND2X2 _14662_ (
    .A(_3827_),
    .B(_3826_),
    .Y(_3804_[11])
);

AND2X2 _14242_ (
    .A(_3607_),
    .B(_3670_),
    .Y(_3606_[0])
);

FILL FILL_1__16169_ (
);

AND2X2 _15867_ (
    .A(_4195__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_4815_)
);

OR2X2 _15447_ (
    .A(_4398_),
    .B(_4401_),
    .Y(_4402_)
);

AND2X2 _15027_ (
    .A(_4008_),
    .B(_4015_),
    .Y(_4016_)
);

OR2X2 _10582_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .B(_1124__bF$buf4),
    .Y(_1100_)
);

FILL FILL_0__10297_ (
);

OR2X2 _10162_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .B(_926__bF$buf1),
    .Y(_880_)
);

FILL FILL_1__17110_ (
);

FILL FILL_1__8719_ (
);

FILL FILL_0__16943_ (
);

FILL FILL_0__16523_ (
);

AND2X2 _19280_ (
    .A(_6255__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_8177_)
);

OR2X2 _8730_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_145_)
);

FILL FILL_1__12089_ (
);

DFFSR _11787_ (
    .CLK(clk_bF$buf51),
    .D(_1653_[9]),
    .Q(\datapath_1.regfile_1.regOut[26] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

OR2X2 _11367_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_1503_)
);

FILL FILL50160x74100 (
);

FILL FILL_1__13450_ (
);

FILL FILL_0__17728_ (
);

FILL FILL_0__17308_ (
);

FILL FILL14440x365560 (
);

FILL FILL199120x39520 (
);

FILL FILL181640x108680 (
);

AND2X2 _9935_ (
    .A(_768_),
    .B(_767_),
    .Y(_729_[19])
);

FILL FILL299440x232180 (
);

AND2X2 _9515_ (
    .A(_548_),
    .B(_547_),
    .Y(_531_[8])
);

FILL FILL18240x286520 (
);

AND2X2 _13933_ (
    .A(_3347__bF$buf2),
    .B(\aluControl_1.inst [2]),
    .Y(_3362_)
);

FILL FILL_0__13648_ (
);

FILL FILL_0__13228_ (
);

OR2X2 _13513_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [8]),
    .Y(_3030_)
);

FILL FILL358720x370500 (
);

FILL FILL386840x103740 (
);

FILL FILL69160x103740 (
);

BUFX2 BUFX2_insert1070 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf4 )
);

BUFX2 BUFX2_insert1071 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf3 )
);

BUFX2 BUFX2_insert1072 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf2 )
);

FILL FILL_0__17061_ (
);

BUFX2 BUFX2_insert1073 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf1 )
);

BUFX2 BUFX2_insert1074 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf0 )
);

BUFX2 BUFX2_insert1075 (
    .A(PCEn),
    .Y(PCEn_bF$buf4)
);

BUFX2 BUFX2_insert1076 (
    .A(PCEn),
    .Y(PCEn_bF$buf3)
);

BUFX2 BUFX2_insert1077 (
    .A(PCEn),
    .Y(PCEn_bF$buf2)
);

BUFX2 BUFX2_insert1078 (
    .A(PCEn),
    .Y(PCEn_bF$buf1)
);

BUFX2 BUFX2_insert1079 (
    .A(PCEn),
    .Y(PCEn_bF$buf0)
);

FILL FILL_1__10155_ (
);

OR2X2 _14718_ (
    .A(\datapath_1.rd1 [30]),
    .B(_3869__bF$buf0),
    .Y(_3865_)
);

FILL FILL86640x113620 (
);

BUFX2 BUFX2_insert890 (
    .A(_3671_),
    .Y(_3671__bF$buf2)
);

BUFX2 BUFX2_insert891 (
    .A(_3671_),
    .Y(_3671__bF$buf1)
);

BUFX2 BUFX2_insert892 (
    .A(_3671_),
    .Y(_3671__bF$buf0)
);

BUFX2 BUFX2_insert893 (
    .A(_6255_),
    .Y(_6255__bF$buf4)
);

FILL FILL_1_CLKBUF1_insert200 (
);

BUFX2 BUFX2_insert894 (
    .A(_6255_),
    .Y(_6255__bF$buf3)
);

FILL FILL_1_CLKBUF1_insert202 (
);

BUFX2 BUFX2_insert895 (
    .A(_6255_),
    .Y(_6255__bF$buf2)
);

BUFX2 BUFX2_insert896 (
    .A(_6255_),
    .Y(_6255__bF$buf1)
);

BUFX2 BUFX2_insert897 (
    .A(_6255_),
    .Y(_6255__bF$buf0)
);

BUFX2 BUFX2_insert898 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf4 )
);

BUFX2 BUFX2_insert899 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf3 )
);

FILL FILL67640x271700 (
);

FILL FILL_0__18686_ (
);

AND2X2 _18971_ (
    .A(_6206__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_7872_)
);

AND2X2 _18551_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_7459_)
);

FILL FILL_0__18266_ (
);

OR2X2 _18131_ (
    .A(_7044_),
    .B(_7043_),
    .Y(_7045_)
);

FILL FILL_0__8787_ (
);

FILL FILL12920x321100 (
);

DFFSR _10638_ (
    .CLK(clk_bF$buf21),
    .D(_1059_[21]),
    .Q(\datapath_1.regfile_1.regOut[17] [21]),
    .R(rst_bF$buf109),
    .S(vdd)
);

OR2X2 _10218_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_917_)
);

OR2X2 _19336_ (
    .A(_8231_),
    .B(_8230_),
    .Y(_8232_)
);

OR2X2 _14891_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [2]),
    .Y(_3940_)
);

DFFSR _14471_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[6]),
    .Q(\datapath_1.Data [6]),
    .R(rst_bF$buf85),
    .S(vdd)
);

AND2X2 _14051_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3463_)
);

FILL FILL60040x4940 (
);

FILL FILL_0__12919_ (
);

FILL FILL_1__16398_ (
);

FILL FILL125400x34580 (
);

FILL FILL141360x286520 (
);

AND2X2 _15676_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_4627_)
);

AND2X2 _15256_ (
    .A(_4213_),
    .B(_4144_),
    .Y(_4214_)
);

OR2X2 _10391_ (
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .Y(_1057_)
);

FILL FILL_0__16332_ (
);

FILL FILL72960x281580 (
);

OR2X2 _11596_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_1652__bF$buf2),
    .Y(_1616_)
);

FILL FILL_1__18544_ (
);

OR2X2 _11176_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .B(_1454__bF$buf3),
    .Y(_1396_)
);

FILL FILL_0__17537_ (
);

AND2X2 _17822_ (
    .A(_6206__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_6741_)
);

AND2X2 _17402_ (
    .A(_6270_),
    .B(\datapath_1.PCJump_27_bF$buf1 ),
    .Y(_6328_)
);

FILL FILL_0__17117_ (
);

FILL FILL_0__12672_ (
);

FILL FILL152000x158080 (
);

FILL FILL_0__12252_ (
);

FILL FILL468920x148200 (
);

DFFSR _9744_ (
    .CLK(clk_bF$buf33),
    .D(_597_[30]),
    .Q(\datapath_1.regfile_1.regOut[10] [30]),
    .R(rst_bF$buf88),
    .S(vdd)
);

OR2X2 _9324_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_461_)
);

FILL FILL129200x34580 (
);

FILL FILL_1__19329_ (
);

FILL FILL468160x375440 (
);

FILL FILL_1__14884_ (
);

FILL FILL_1__14464_ (
);

OR2X2 _18607_ (
    .A(_7513_),
    .B(_7512_),
    .Y(_7514_)
);

FILL FILL299440x370500 (
);

FILL FILL_0__13877_ (
);

FILL FILL_0__13457_ (
);

AND2X2 _13742_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3216_)
);

AND2X2 _13322_ (
    .A(_2862_),
    .B(_2204_),
    .Y(_2863_)
);

FILL FILL438520x29640 (
);

FILL FILL208240x247000 (
);

FILL FILL_0__17290_ (
);

FILL FILL_1__15249_ (
);

FILL FILL57000x163020 (
);

AND2X2 _14947_ (
    .A(_3977_),
    .B(_3976_),
    .Y(_3936_[20])
);

AND2X2 _14527_ (
    .A(_3757_),
    .B(_3756_),
    .Y(_3738_[9])
);

AND2X2 _14107_ (
    .A(_3344__bF$buf1),
    .B(gnd),
    .Y(_3511_)
);

FILL FILL160360x34580 (
);

FILL FILL259160x9880 (
);

FILL FILL_1__16610_ (
);

FILL FILL_1__19082_ (
);

AND2X2 _18780_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_7684_)
);

FILL FILL_0__18495_ (
);

AND2X2 _18360_ (
    .A(_6328__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_7271_)
);

FILL FILL431680x103740 (
);

FILL FILL267520x19760 (
);

FILL FILL_0__8596_ (
);

OR2X2 _10867_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_1256__bF$buf2),
    .Y(_1250_)
);

OR2X2 _10447_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .B(_1058__bF$buf1),
    .Y(_1030_)
);

OR2X2 _10027_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .B(_860__bF$buf3),
    .Y(_810_)
);

FILL FILL_1__12950_ (
);

FILL FILL_0__16808_ (
);

FILL FILL_0__11943_ (
);

OR2X2 _19145_ (
    .A(_8036_),
    .B(_8043_),
    .Y(_8044_)
);

OR2X2 _14280_ (
    .A(\datapath_1.ALUResult [13]),
    .B(_3671__bF$buf3),
    .Y(_3633_)
);

FILL FILL_1__13315_ (
);

FILL FILL260680x172900 (
);

OR2X2 _15485_ (
    .A(_4437_),
    .B(_4438_),
    .Y(_4439_)
);

AND2X2 _15065_ (
    .A(_4053_),
    .B(_4029_),
    .Y(\datapath_1.regfile_1.regEn [1])
);

FILL FILL_0__16981_ (
);

FILL FILL_0__16561_ (
);

FILL FILL_0__16141_ (
);

FILL FILL225720x49400 (
);

FILL FILL_0__17766_ (
);

AND2X2 _17631_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_6553_)
);

AND2X2 _17211_ (
    .A(_4236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_6138_)
);

FILL FILL249280x153140 (
);

FILL FILL262200x340860 (
);

DFFSR _9973_ (
    .CLK(clk_bF$buf1),
    .D(_729_[1]),
    .Q(\datapath_1.regfile_1.regOut[12] [1]),
    .R(rst_bF$buf96),
    .S(vdd)
);

OR2X2 _9553_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .B(_596__bF$buf0),
    .Y(_574_)
);

OR2X2 _9133_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .B(_398__bF$buf3),
    .Y(_354_)
);

FILL FILL_1__14273_ (
);

OR2X2 _18836_ (
    .A(_7732_),
    .B(_7739_),
    .Y(_7740_)
);

FILL FILL_0_BUFX2_insert531 (
);

AND2X2 _18416_ (
    .A(_6244__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_7326_)
);

FILL FILL_0_BUFX2_insert533 (
);

AND2X2 _13971_ (
    .A(_3352__bF$buf0),
    .B(\aluControl_1.inst [5]),
    .Y(_3395_)
);

FILL FILL_0__13266_ (
);

FILL FILL_0_BUFX2_insert535 (
);

AND2X2 _13551_ (
    .A(_3055_),
    .B(_3054_),
    .Y(_1_[20])
);

FILL FILL_0_BUFX2_insert536 (
);

AND2X2 _13131_ (
    .A(_2683_),
    .B(_2671_),
    .Y(_2684_)
);

FILL FILL_0_BUFX2_insert537 (
);

FILL FILL_0_BUFX2_insert538 (
);

FILL FILL_0_BUFX2_insert539 (
);

FILL FILL229520x49400 (
);

FILL FILL397480x44460 (
);

FILL FILL_1__15898_ (
);

INVX2 _14756_ (
    .A(vdd),
    .Y(_3935_)
);

DFFSR _14336_ (
    .CLK(clk_bF$buf62),
    .D(_3606_[0]),
    .Q(ALUOut[0]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL484880x153140 (
);

FILL FILL220400x202540 (
);

FILL FILL_0__15832_ (
);

FILL FILL_0__15412_ (
);

FILL FILL126160x64220 (
);

FILL FILL439280x276640 (
);

FILL FILL97280x158080 (
);

AND2X2 _10676_ (
    .A(_1142_),
    .B(_1141_),
    .Y(_1125_[8])
);

DFFSR _10256_ (
    .CLK(clk_bF$buf54),
    .D(_861_[26]),
    .Q(\datapath_1.regfile_1.regOut[14] [26]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL_0__16617_ (
);

AND2X2 _16902_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_5834_)
);

FILL FILL_0__11752_ (
);

OR2X2 _19374_ (
    .A(_8268_),
    .B(_8265_),
    .Y(_8269_)
);

FILL FILL_0__19089_ (
);

FILL FILL114760x340860 (
);

DFFSR _8824_ (
    .CLK(clk_bF$buf61),
    .D(_135_[13]),
    .Q(\datapath_1.regfile_1.regOut[3] [13]),
    .R(rst_bF$buf55),
    .S(vdd)
);

BUFX2 _8404_ (
    .A(_1_[12]),
    .Y(memoryAddress[12])
);

FILL FILL38000x202540 (
);

FILL FILL120080x88920 (
);

FILL FILL_1__18409_ (
);

FILL FILL182400x69160 (
);

FILL FILL502360x98800 (
);

FILL FILL_0__12957_ (
);

NAND3X1 _12822_ (
    .A(_2386_),
    .B(ALUControl[1]),
    .C(_2154_),
    .Y(_2387_)
);

FILL FILL_0__12537_ (
);

OR2X2 _12402_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_2033_)
);

FILL FILL_0__12117_ (
);

FILL FILL15960x103740 (
);

AND2X2 _15294_ (
    .A(_4187__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_4251_)
);

DFFSR _9609_ (
    .CLK(clk_bF$buf97),
    .D(_531_[24]),
    .Q(\datapath_1.regfile_1.regOut[9] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL_0__16790_ (
);

FILL FILL_0__16370_ (
);

OR2X2 _13607_ (
    .A(_3098_),
    .B(_3099_),
    .Y(_3100_)
);

AND2X2 _16499_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_5438_)
);

OR2X2 _16079_ (
    .A(_5022_),
    .B(_5023_),
    .Y(_5024_)
);

FILL FILL_1__18582_ (
);

FILL FILL_1__18162_ (
);

OR2X2 _17860_ (
    .A(_6775_),
    .B(_6778_),
    .Y(_6779_)
);

FILL FILL281960x222300 (
);

OR2X2 _17440_ (
    .A(_6364_),
    .B(_6350_),
    .Y(_6365_)
);

FILL FILL_0__17155_ (
);

AND2X2 _17020_ (
    .A(_4160__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_5950_)
);

FILL FILL440040x187720 (
);

FILL FILL_0__12290_ (
);

AND2X2 _9782_ (
    .A(_686_),
    .B(_685_),
    .Y(_663_[11])
);

AND2X2 _9362_ (
    .A(_466_),
    .B(_529_),
    .Y(_465_[0])
);

FILL FILL454480x148200 (
);

AND2X2 _18645_ (
    .A(_7551_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd1 [19])
);

FILL FILL490960x321100 (
);

AND2X2 _18225_ (
    .A(_6232__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_7138_)
);

FILL FILL_0__13495_ (
);

AND2X2 _13780_ (
    .A(_3081__bF$buf1),
    .B(ALUOut[27]),
    .Y(_3248_)
);

NAND2X1 _13360_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2899_)
);

FILL FILL_0__19301_ (
);

FILL FILL_1__12815_ (
);

FILL FILL_0__9822_ (
);

FILL FILL_0__9402_ (
);

FILL FILL_1__15287_ (
);

FILL FILL328320x281580 (
);

DFFSR _14985_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[4]),
    .Q(\datapath_1.mux_iord.din0 [4]),
    .R(rst_bF$buf18),
    .S(vdd)
);

OR2X2 _14565_ (
    .A(memoryOutData[22]),
    .B(_3803__bF$buf3),
    .Y(_3783_)
);

AND2X2 _14145_ (
    .A(_3541_),
    .B(_3604_),
    .Y(\datapath_1.mux_wd3.dout [0])
);

FILL FILL110960x370500 (
);

FILL FILL_0__15641_ (
);

FILL FILL133000x335920 (
);

FILL FILL488680x167960 (
);

FILL FILL247760x202540 (
);

OR2X2 _10485_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_1055_)
);

OR2X2 _10065_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_835_)
);

FILL FILL_0__16846_ (
);

OR2X2 _16711_ (
    .A(_5644_),
    .B(_5645_),
    .Y(_5646_)
);

FILL FILL_0__16006_ (
);

FILL FILL_0__11981_ (
);

AND2X2 _19183_ (
    .A(_6321__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_8081_)
);

FILL FILL414960x375440 (
);

AND2X2 _8633_ (
    .A(_100_),
    .B(_99_),
    .Y(_69_[15])
);

FILL FILL372400x49400 (
);

FILL FILL_1__13773_ (
);

AND2X2 _17916_ (
    .A(_6302__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_6834_)
);

FILL FILL_0__12766_ (
);

XOR2X1 _12631_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2196_)
);

FILL FILL_0__12346_ (
);

OR2X2 _12211_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .B(_1982__bF$buf4),
    .Y(_1926_)
);

FILL FILL121600x108680 (
);

FILL FILL7600x261820 (
);

OR2X2 _9838_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_728__bF$buf1),
    .Y(_724_)
);

OR2X2 _9418_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_530__bF$buf4),
    .Y(_504_)
);

FILL FILL_1__14138_ (
);

AND2X2 _13836_ (
    .A(_3290_),
    .B(_3289_),
    .Y(\datapath_1.alu_1.ALUInA [6])
);

OR2X2 _13416_ (
    .A(_2389_),
    .B(_2376__bF$buf1),
    .Y(_2951_)
);

FILL FILL467400x74100 (
);

FILL FILL_0__14912_ (
);

FILL FILL104880x79040 (
);

FILL FILL76760x365560 (
);

FILL FILL343520x153140 (
);

FILL FILL_0__17384_ (
);

FILL FILL_1__10058_ (
);

FILL FILL243200x247000 (
);

FILL FILL_1__16704_ (
);

DFFSR _9591_ (
    .CLK(clk_bF$buf29),
    .D(_531_[6]),
    .Q(\datapath_1.regfile_1.regOut[9] [6]),
    .R(rst_bF$buf40),
    .S(vdd)
);

OR2X2 _9171_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_379_)
);

FILL FILL_0__10832_ (
);

AND2X2 _18874_ (
    .A(_6255__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_7777_)
);

FILL FILL_0__18589_ (
);

FILL FILL_0__18169_ (
);

FILL FILL_0_BUFX2_insert911 (
);

AND2X2 _18454_ (
    .A(_6287__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_7363_)
);

AND2X2 _18034_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_6950_)
);

FILL FILL_0_BUFX2_insert913 (
);

FILL FILL_0_BUFX2_insert915 (
);

FILL FILL_0_BUFX2_insert916 (
);

FILL FILL_0_BUFX2_insert917 (
);

FILL FILL17480x217360 (
);

FILL FILL_0_BUFX2_insert918 (
);

FILL FILL_0_BUFX2_insert919 (
);

FILL FILL_1__17909_ (
);

FILL FILL_0__9631_ (
);

OR2X2 _11902_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .B(_1784__bF$buf1),
    .Y(_1780_)
);

AND2X2 _19239_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_8136_)
);

FILL FILL338960x138320 (
);

AND2X2 _14794_ (
    .A(_3895_),
    .B(_3894_),
    .Y(_3870_[12])
);

FILL FILL_0__14089_ (
);

AND2X2 _14374_ (
    .A(_3675_),
    .B(_3674_),
    .Y(_3672_[1])
);

FILL FILL_0__15450_ (
);

FILL FILL_0__15030_ (
);

FILL FILL374680x217360 (
);

FILL FILL427880x54340 (
);

FILL FILL364040x177840 (
);

AND2X2 _15999_ (
    .A(_4223__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_4945_)
);

AND2X2 _15579_ (
    .A(_4228__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_4532_)
);

NOR2X1 _15159_ (
    .A(_4042_),
    .B(_4005_),
    .Y(_4122_)
);

FILL FILL_1__17662_ (
);

OR2X2 _10294_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .B(_992__bF$buf3),
    .Y(_948_)
);

FILL FILL_0__16655_ (
);

AND2X2 _16940_ (
    .A(_4195__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_5872_)
);

OR2X2 _16520_ (
    .A(_5457_),
    .B(_5454_),
    .Y(_5458_)
);

FILL FILL_0__16235_ (
);

AND2X2 _16100_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_5045_)
);

FILL FILL_0__11370_ (
);

FILL FILL23560x79040 (
);

FILL FILL104120x370500 (
);

FILL FILL134520x281580 (
);

FILL FILL112480x83980 (
);

OR2X2 _8862_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_213_)
);

BUFX2 _8442_ (
    .A(_2_[18]),
    .Y(memoryWriteData[18])
);

FILL FILL177840x345800 (
);

OR2X2 _11499_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_1571_)
);

OR2X2 _11079_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_1351_)
);

FILL FILL_1__18027_ (
);

AND2X2 _17725_ (
    .A(_6300__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_6646_)
);

AND2X2 _17305_ (
    .A(_6226_),
    .B(_6204_),
    .Y(_6231_)
);

FILL FILL_0__12995_ (
);

AND2X2 _12860_ (
    .A(_2423_),
    .B(_2424_),
    .Y(_2425_)
);

DFFSR _12440_ (
    .CLK(clk_bF$buf15),
    .D(_1983_[17]),
    .Q(\datapath_1.regfile_1.regOut[31] [17]),
    .R(rst_bF$buf31),
    .S(vdd)
);

AND2X2 _12020_ (
    .A(_1838_),
    .B(_1837_),
    .Y(_1785_[26])
);

FILL FILL_0__18801_ (
);

FILL FILL276640x59280 (
);

AND2X2 _9647_ (
    .A(_616_),
    .B(_615_),
    .Y(_597_[9])
);

DFFSR _9227_ (
    .CLK(clk_bF$buf53),
    .D(_333_[29]),
    .Q(\datapath_1.regfile_1.regOut[6] [29]),
    .R(rst_bF$buf111),
    .S(vdd)
);

FILL FILL_0__8902_ (
);

FILL FILL212800x79040 (
);

OR2X2 _13645_ (
    .A(_3132_),
    .B(_3131_),
    .Y(_3133_)
);

NOR3X1 _13225_ (
    .A(_2768_),
    .B(_2769_),
    .C(_2771_),
    .Y(_2772_)
);

FILL FILL27360x79040 (
);

FILL FILL116280x83980 (
);

FILL FILL13680x247000 (
);

FILL FILL129960x266760 (
);

FILL FILL_0__14301_ (
);

FILL FILL330600x345800 (
);

FILL FILL266760x326040 (
);

FILL FILL153520x4940 (
);

FILL FILL_0_CLKBUF1_insert141 (
);

FILL FILL_0__15926_ (
);

FILL FILL_0__15506_ (
);

FILL FILL_0_CLKBUF1_insert143 (
);

FILL FILL_0_CLKBUF1_insert144 (
);

FILL FILL_0_CLKBUF1_insert145 (
);

FILL FILL440800x29640 (
);

FILL FILL_0_CLKBUF1_insert146 (
);

FILL FILL_0_CLKBUF1_insert147 (
);

FILL FILL_0_CLKBUF1_insert148 (
);

FILL FILL_0__10221_ (
);

FILL FILL210520x0 (
);

OR2X2 _18683_ (
    .A(_7588_),
    .B(_7585_),
    .Y(_7589_)
);

AND2X2 _18263_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_7175_)
);

FILL FILL233320x29640 (
);

FILL FILL10640x143260 (
);

FILL FILL408120x39520 (
);

FILL FILL_0__9440_ (
);

AND2X2 _11711_ (
    .A(_1672_),
    .B(_1671_),
    .Y(_1653_[9])
);

FILL FILL_0__11426_ (
);

FILL FILL_0__9020_ (
);

AND2X2 _19468_ (
    .A(_8347_),
    .B(_8346_),
    .Y(_8320_[13])
);

AND2X2 _19048_ (
    .A(_6323__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_7948_)
);

OR2X2 _14183_ (
    .A(\datapath_1.Data [13]),
    .B(_3605__bF$buf3),
    .Y(_3567_)
);

AND2X2 _8918_ (
    .A(_250_),
    .B(_249_),
    .Y(_201_[24])
);

FILL FILL214320x148200 (
);

FILL FILL305520x350740 (
);

FILL FILL_1__13638_ (
);

FILL FILL478040x197600 (
);

FILL FILL_1_BUFX2_insert460 (
);

OAI21X1 _12916_ (
    .A(_2331_),
    .B(_2329_),
    .C(_2327_),
    .Y(_2481_)
);

FILL FILL_1_BUFX2_insert468 (
);

FILL FILL250040x227240 (
);

OR2X2 _15388_ (
    .A(_4343_),
    .B(_4342_),
    .Y(_4344_)
);

FILL FILL_1__17051_ (
);

FILL FILL_0__16884_ (
);

FILL FILL497040x0 (
);

FILL FILL153520x261820 (
);

OR2X2 _8671_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .B(_134__bF$buf1),
    .Y(_126_)
);

FILL FILL31920x261820 (
);

FILL FILL_1__18676_ (
);

FILL FILL_1__13391_ (
);

FILL FILL_0__17669_ (
);

AND2X2 _17954_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_6871_)
);

FILL FILL_0__17249_ (
);

OR2X2 _17534_ (
    .A(_6457_),
    .B(_6456_),
    .Y(_6458_)
);

AND2X2 _17114_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_6043_)
);

FILL FILL31160x167960 (
);

FILL FILL_0__18610_ (
);

INVX2 _9876_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .Y(_794_)
);

DFFSR _9456_ (
    .CLK(clk_bF$buf99),
    .D(_465_[0]),
    .Q(\datapath_1.regfile_1.regOut[8] [0]),
    .R(rst_bF$buf19),
    .S(vdd)
);

OR2X2 _9036_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_309_)
);

OR2X2 _18739_ (
    .A(_7643_),
    .B(_7636_),
    .Y(_7644_)
);

OR2X2 _18319_ (
    .A(_7197_),
    .B(_7230_),
    .Y(_7231_)
);

OR2X2 _13874_ (
    .A(\datapath_1.a [19]),
    .B(_3342__bF$buf3),
    .Y(_3316_)
);

FILL FILL_0__13589_ (
);

AND2X2 _13454_ (
    .A(_2963_),
    .B(_2973_),
    .Y(_2987_)
);

FILL FILL216600x301340 (
);

FILL FILL105640x182780 (
);

INVX1 _13034_ (
    .A(_2331_),
    .Y(_2592_)
);

FILL FILL_0__14110_ (
);

FILL FILL242440x242060 (
);

FILL FILL279680x365560 (
);

FILL FILL_1__10096_ (
);

AND2X2 _14659_ (
    .A(_3825_),
    .B(_3824_),
    .Y(_3804_[10])
);

OR2X2 _14239_ (
    .A(ALUOut[0]),
    .B(vdd),
    .Y(_3670_)
);

FILL FILL_0__15735_ (
);

FILL FILL_0__15315_ (
);

AND2X2 _15600_ (
    .A(_4142__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [5]),
    .Y(_4553_)
);

FILL FILL_0__10870_ (
);

FILL FILL_0__10450_ (
);

FILL FILL_0__10030_ (
);

AND2X2 _18492_ (
    .A(_6244__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_7401_)
);

AND2X2 _18072_ (
    .A(_6321__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_6987_)
);

FILL FILL430160x93860 (
);

OR2X2 _10999_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .B(_1322__bF$buf4),
    .Y(_1318_)
);

FILL FILL_1__17527_ (
);

OR2X2 _10579_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .B(_1124__bF$buf1),
    .Y(_1098_)
);

OR2X2 _10159_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .B(_926__bF$buf4),
    .Y(_878_)
);

AND2X2 _16805_ (
    .A(_4210__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_5739_)
);

INVX2 _11940_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .Y(_1850_)
);

FILL FILL_0__11235_ (
);

DFFSR _11520_ (
    .CLK(clk_bF$buf99),
    .D(_1521_[0]),
    .Q(\datapath_1.regfile_1.regOut[24] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

OR2X2 _11100_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_1365_)
);

AND2X2 _19277_ (
    .A(_6259__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_8174_)
);

FILL FILL282720x202540 (
);

OR2X2 _8727_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_143_)
);

FILL FILL432440x365560 (
);

FILL FILL_1__13867_ (
);

INVX1 _12725_ (
    .A(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2290_)
);

DFFSR _12305_ (
    .CLK(clk_bF$buf45),
    .D(_1917_[11]),
    .Q(\datapath_1.regfile_1.regOut[30] [11]),
    .R(rst_bF$buf54),
    .S(vdd)
);

AND2X2 _15197_ (
    .A(_4154__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_4155_)
);

FILL FILL_0__13801_ (
);

FILL FILL_1__17280_ (
);

FILL FILL436240x286520 (
);

FILL FILL_1__8469_ (
);

FILL FILL_0__16273_ (
);

FILL FILL_1__9830_ (
);

AND2X2 _8480_ (
    .A(_18_),
    .B(_17_),
    .Y(_3_[7])
);

FILL FILL113240x98800 (
);

FILL FILL286520x83980 (
);

FILL FILL_0__17898_ (
);

FILL FILL_0__17478_ (
);

OR2X2 _17763_ (
    .A(_6682_),
    .B(_6679_),
    .Y(_6683_)
);

OR2X2 _17343_ (
    .A(_6268_),
    .B(_6242_),
    .Y(_6269_)
);

FILL FILL206720x256880 (
);

OR2X2 _9685_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .B(_662__bF$buf0),
    .Y(_642_)
);

OR2X2 _9265_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_464__bF$buf3),
    .Y(_422_)
);

FILL FILL_1_CLKBUF1_insert174 (
);

FILL FILL_1_CLKBUF1_insert176 (
);

FILL FILL_1_CLKBUF1_insert178 (
);

FILL FILL_0__8520_ (
);

FILL FILL_0__10926_ (
);

OR2X2 _18968_ (
    .A(_7837_),
    .B(_7869_),
    .Y(_7870_)
);

AND2X2 _18548_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_7456_)
);

OR2X2 _18128_ (
    .A(_7041_),
    .B(_7040_),
    .Y(_7042_)
);

FILL FILL_0__13398_ (
);

AND2X2 _13683_ (
    .A(_3084__bF$buf4),
    .B(\datapath_1.PCJump [13]),
    .Y(_3165_)
);

INVX1 _13263_ (
    .A(_2807_),
    .Y(\datapath_1.ALUResult [11])
);

FILL FILL_0__9305_ (
);

OR2X2 _14888_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [1]),
    .Y(_3938_)
);

DFFSR _14468_ (
    .CLK(clk_bF$buf2),
    .D(_3672_[3]),
    .Q(\datapath_1.Data [3]),
    .R(rst_bF$buf26),
    .S(vdd)
);

AND2X2 _14048_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3461_)
);

FILL FILL_1__16131_ (
);

FILL FILL_0__15964_ (
);

FILL FILL_0__15124_ (
);

FILL FILL428640x167960 (
);

FILL FILL92720x311220 (
);

DFFSR _10388_ (
    .CLK(clk_bF$buf0),
    .D(_927_[29]),
    .Q(\datapath_1.regfile_1.regOut[15] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

FILL FILL_1__12891_ (
);

FILL FILL475000x54340 (
);

FILL FILL_0__16749_ (
);

OR2X2 _16614_ (
    .A(_5549_),
    .B(_5550_),
    .Y(_5551_)
);

FILL FILL_0__16329_ (
);

FILL FILL_0__11884_ (
);

FILL FILL_0__11044_ (
);

AND2X2 _19086_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_7986_)
);

DFFSR _8956_ (
    .CLK(clk_bF$buf64),
    .D(_201_[16]),
    .Q(\datapath_1.regfile_1.regOut[4] [16]),
    .R(rst_bF$buf10),
    .S(vdd)
);

OR2X2 _8536_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .B(_68__bF$buf3),
    .Y(_56_)
);

FILL FILL_1__13256_ (
);

AND2X2 _17819_ (
    .A(_6211__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_6738_)
);

FILL FILL130720x247000 (
);

OAI21X1 _12954_ (
    .A(_2354_),
    .B(_2376__bF$buf3),
    .C(_2516_),
    .Y(_2517_)
);

FILL FILL_0__12249_ (
);

AND2X2 _12534_ (
    .A(_2123_),
    .B(_2118_),
    .Y(_2124_)
);

OR2X2 _12114_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_1881_)
);

FILL FILL_1_BUFX2_insert848 (
);

FILL FILL_0__16082_ (
);

FILL FILL422560x108680 (
);

AND2X2 _13739_ (
    .A(_3084__bF$buf0),
    .B(\datapath_1.PCJump [21]),
    .Y(_3213_)
);

NAND3X1 _13319_ (
    .A(_2859_),
    .B(_2189_),
    .C(_2190_),
    .Y(_2860_)
);

FILL FILL_1__15822_ (
);

FILL FILL253840x103740 (
);

FILL FILL48640x153140 (
);

FILL FILL18240x69160 (
);

FILL FILL_0__14815_ (
);

BUFX2 BUFX2_insert510 (
    .A(_4195_),
    .Y(_4195__bF$buf0)
);

BUFX2 BUFX2_insert511 (
    .A(_6206_),
    .Y(_6206__bF$buf4)
);

BUFX2 BUFX2_insert512 (
    .A(_6206_),
    .Y(_6206__bF$buf3)
);

BUFX2 BUFX2_insert513 (
    .A(_6206_),
    .Y(_6206__bF$buf2)
);

OR2X2 _17992_ (
    .A(_6908_),
    .B(_6892_),
    .Y(_6909_)
);

BUFX2 BUFX2_insert514 (
    .A(_6206_),
    .Y(_6206__bF$buf1)
);

AND2X2 _17572_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_6495_)
);

BUFX2 BUFX2_insert515 (
    .A(_6206_),
    .Y(_6206__bF$buf0)
);

FILL FILL_0__17287_ (
);

BUFX2 BUFX2_insert516 (
    .A(_3084_),
    .Y(_3084__bF$buf4)
);

OR2X2 _17152_ (
    .A(_6079_),
    .B(_6078_),
    .Y(_6080_)
);

BUFX2 BUFX2_insert517 (
    .A(_3084_),
    .Y(_3084__bF$buf3)
);

BUFX2 BUFX2_insert518 (
    .A(_3084_),
    .Y(_3084__bF$buf2)
);

BUFX2 BUFX2_insert519 (
    .A(_3084_),
    .Y(_3084__bF$buf1)
);

FILL FILL386840x98800 (
);

FILL FILL234080x167960 (
);

AND2X2 _9494_ (
    .A(_534_),
    .B(_533_),
    .Y(_531_[1])
);

DFFSR _9074_ (
    .CLK(clk_bF$buf59),
    .D(_267_[5]),
    .Q(\datapath_1.regfile_1.regOut[5] [5]),
    .R(rst_bF$buf106),
    .S(vdd)
);

FILL FILL_1__19499_ (
);

OR2X2 _10600_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_1124__bF$buf3),
    .Y(_1112_)
);

FILL FILL_0__10315_ (
);

FILL FILL_0_BUFX2_insert31 (
);

AND2X2 _18777_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_7681_)
);

OR2X2 _18357_ (
    .A(_7267_),
    .B(_7266_),
    .Y(_7268_)
);

FILL FILL_0_BUFX2_insert33 (
);

FILL FILL_0_BUFX2_insert34 (
);

FILL FILL_0_BUFX2_insert35 (
);

FILL FILL_0_BUFX2_insert36 (
);

FILL FILL_0_BUFX2_insert37 (
);

OR2X2 _13492_ (
    .A(IorD_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [1]),
    .Y(_3016_)
);

NAND2X1 _13072_ (
    .A(_2264_),
    .B(_2504_),
    .Y(_2628_)
);

FILL FILL_0_BUFX2_insert39 (
);

FILL FILL_0__19433_ (
);

FILL FILL_0__19013_ (
);

FILL FILL_1__12527_ (
);

FILL FILL_0__9954_ (
);

FILL FILL_0__9534_ (
);

FILL FILL_0__9114_ (
);

DFFSR _11805_ (
    .CLK(clk_bF$buf70),
    .D(_1653_[27]),
    .Q(\datapath_1.regfile_1.regOut[26] [27]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL88920x113620 (
);

OR2X2 _14697_ (
    .A(\datapath_1.rd1 [23]),
    .B(_3869__bF$buf2),
    .Y(_3851_)
);

OR2X2 _14277_ (
    .A(\datapath_1.ALUResult [12]),
    .B(_3671__bF$buf2),
    .Y(_3631_)
);

FILL FILL291840x271700 (
);

FILL FILL_1__16780_ (
);

FILL FILL369360x167960 (
);

FILL FILL_0__15773_ (
);

FILL FILL_0__15353_ (
);

FILL FILL_1__8910_ (
);

FILL FILL209760x64220 (
);

OR2X2 _10197_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_903_)
);

FILL FILL_1__17145_ (
);

FILL FILL_1__12280_ (
);

FILL FILL_0__16978_ (
);

FILL FILL14440x227240 (
);

AND2X2 _16843_ (
    .A(_4175__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_5776_)
);

FILL FILL_0__16138_ (
);

OR2X2 _16423_ (
    .A(_5359_),
    .B(_5362_),
    .Y(_5363_)
);

AND2X2 _16003_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_4949_)
);

FILL FILL_0__11693_ (
);

AND2X2 _8765_ (
    .A(_168_),
    .B(_167_),
    .Y(_135_[16])
);

FILL FILL148200x34580 (
);

AND2X2 _17628_ (
    .A(_6206__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_6550_)
);

OR2X2 _17208_ (
    .A(_6120_),
    .B(_6135_),
    .Y(_6136_)
);

FILL FILL143640x286520 (
);

INVX1 _12763_ (
    .A(_2327_),
    .Y(_2328_)
);

FILL FILL_0__12478_ (
);

OR2X2 _12343_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .B(_2048__bF$buf1),
    .Y(_1994_)
);

FILL FILL437760x14820 (
);

FILL FILL_0__8805_ (
);

FILL FILL380760x118560 (
);

AND2X2 _13968_ (
    .A(_3347__bF$buf0),
    .B(\datapath_1.PCJump [9]),
    .Y(_3392_)
);

AND2X2 _13548_ (
    .A(_3053_),
    .B(_3052_),
    .Y(_1_[19])
);

AND2X2 _13128_ (
    .A(_2680_),
    .B(_2676_),
    .Y(_2681_)
);

FILL FILL_0__14204_ (
);

INVX1 _17381_ (
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_6307_)
);

FILL FILL_0__17096_ (
);

FILL FILL206720x326040 (
);

FILL FILL61560x286520 (
);

FILL FILL213560x9880 (
);

FILL FILL207480x88920 (
);

FILL FILL_1__11971_ (
);

FILL FILL_0__15829_ (
);

FILL FILL_0__10964_ (
);

FILL FILL375440x335920 (
);

OR2X2 _18586_ (
    .A(_7492_),
    .B(_7491_),
    .Y(_7493_)
);

AND2X2 _18166_ (
    .A(_6221__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_7080_)
);

FILL FILL316160x321100 (
);

FILL FILL_0__19242_ (
);

FILL FILL232560x9880 (
);

FILL FILL_1__12756_ (
);

FILL FILL_1__12336_ (
);

FILL FILL_0__9763_ (
);

FILL FILL395200x232180 (
);

OR2X2 _11614_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .B(_1652__bF$buf3),
    .Y(_1628_)
);

FILL FILL_0__11329_ (
);

FILL FILL456000x202540 (
);

AND2X2 _14086_ (
    .A(_3344__bF$buf1),
    .B(gnd),
    .Y(_3493_)
);

FILL FILL428640x237120 (
);

AND2X2 _12819_ (
    .A(_2383_),
    .B(_2158_),
    .Y(_2384_)
);

FILL FILL72960x143260 (
);

FILL FILL158840x251940 (
);

FILL FILL_1__17794_ (
);

FILL FILL_0__16787_ (
);

OR2X2 _16652_ (
    .A(_5586_),
    .B(_5587_),
    .Y(_5588_)
);

FILL FILL_0__16367_ (
);

OR2X2 _16232_ (
    .A(_5167_),
    .B(_5174_),
    .Y(_5175_)
);

FILL FILL_0__11082_ (
);

FILL FILL_1__9924_ (
);

OR2X2 _8994_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_281_)
);

DFFSR _8574_ (
    .CLK(clk_bF$buf34),
    .D(_3_[21]),
    .Q(\datapath_1.regfile_1.regOut[1] [21]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_1__18999_ (
);

AND2X2 _17857_ (
    .A(_6300__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_6776_)
);

OR2X2 _17437_ (
    .A(_6361_),
    .B(_6360_),
    .Y(_6362_)
);

FILL FILL253840x4940 (
);

OR2X2 _17017_ (
    .A(_5947_),
    .B(_5916_),
    .Y(_5948_)
);

INVX1 _12992_ (
    .A(_2481_),
    .Y(_2553_)
);

INVX1 _12572_ (
    .A(vdd),
    .Y(_2145_)
);

FILL FILL_0__12287_ (
);

AND2X2 _12152_ (
    .A(_1906_),
    .B(_1905_),
    .Y(_1851_[27])
);

FILL FILL_0__18933_ (
);

FILL FILL_0__18513_ (
);

AND2X2 _9779_ (
    .A(_684_),
    .B(_683_),
    .Y(_663_[10])
);

FILL FILL76760x251940 (
);

OR2X2 _9359_ (
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .Y(_529_)
);

FILL FILL_1__11607_ (
);

FILL FILL_1__14079_ (
);

AND2X2 _13777_ (
    .A(_3089__bF$buf0),
    .B(gnd),
    .Y(_3246_)
);

NAND3X1 _13357_ (
    .A(ALUControl[1]),
    .B(\datapath_1.alu_1.ALUInB [5]),
    .C(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2896_)
);

FILL FILL_0__14433_ (
);

OR2X2 _17190_ (
    .A(_6117_),
    .B(_6116_),
    .Y(_6118_)
);

FILL FILL_1__16645_ (
);

FILL FILL_1__11360_ (
);

FILL FILL306280x276640 (
);

FILL FILL281960x158080 (
);

AND2X2 _15923_ (
    .A(_4146__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_4871_)
);

OR2X2 _15503_ (
    .A(_4456_),
    .B(_4455_),
    .Y(_4457_)
);

FILL FILL_0__15218_ (
);

FILL FILL51680x163020 (
);

OR2X2 _18395_ (
    .A(_7303_),
    .B(_7304_),
    .Y(_7305_)
);

FILL FILL_0__19051_ (
);

FILL FILL_1__12985_ (
);

OR2X2 _16708_ (
    .A(_5641_),
    .B(_5642_),
    .Y(_5643_)
);

FILL FILL_0__11978_ (
);

FILL FILL_0__9572_ (
);

FILL FILL_0__11558_ (
);

FILL FILL_0__9152_ (
);

AND2X2 _11843_ (
    .A(_1740_),
    .B(_1739_),
    .Y(_1719_[10])
);

OR2X2 _11423_ (
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .Y(_1585_)
);

AND2X2 _11003_ (
    .A(_1320_),
    .B(_1319_),
    .Y(_1257_[31])
);

FILL FILL373160x14820 (
);

FILL FILL86640x93860 (
);

FILL FILL_0__15391_ (
);

OR2X2 _12628_ (
    .A(_2192_),
    .B(_2185_),
    .Y(_2193_)
);

FILL FILL300960x311220 (
);

OR2X2 _12208_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .B(_1982__bF$buf4),
    .Y(_1924_)
);

FILL FILL91960x123500 (
);

FILL FILL_0__13704_ (
);

FILL FILL_0__16596_ (
);

AND2X2 _16881_ (
    .A(_4177__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_5814_)
);

FILL FILL_0__16176_ (
);

AND2X2 _16461_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_5400_)
);

AND2X2 _16041_ (
    .A(_4158__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_4987_)
);

OR2X2 _17666_ (
    .A(_6580_),
    .B(_6587_),
    .Y(_6588_)
);

FILL FILL34200x355680 (
);

AND2X2 _17246_ (
    .A(_4225__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_6173_)
);

OR2X2 _12381_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_2019_)
);

FILL FILL_0__12096_ (
);

DFFSR _9588_ (
    .CLK(clk_bF$buf27),
    .D(_531_[3]),
    .Q(\datapath_1.regfile_1.regOut[9] [3]),
    .R(rst_bF$buf28),
    .S(vdd)
);

FILL FILL17480x330980 (
);

OR2X2 _9168_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_377_)
);

FILL FILL235600x9880 (
);

FILL FILL_0__8843_ (
);

FILL FILL_0__10829_ (
);

FILL FILL_0__10409_ (
);

FILL FILL_0_BUFX2_insert880 (
);

FILL FILL_0_BUFX2_insert881 (
);

FILL FILL_0_BUFX2_insert882 (
);

FILL FILL_0_BUFX2_insert884 (
);

AND2X2 _13586_ (
    .A(_3080_),
    .B(ALUOp[0]),
    .Y(_3081_)
);

FILL FILL_0_BUFX2_insert886 (
);

OR2X2 _13166_ (
    .A(_2157__bF$buf2),
    .B(_2715_),
    .Y(_2716_)
);

FILL FILL_0_BUFX2_insert888 (
);

FILL FILL_0__19107_ (
);

FILL FILL442320x187720 (
);

FILL FILL_0__14242_ (
);

FILL FILL283480x128440 (
);

FILL FILL_0__15867_ (
);

FILL FILL_0__15447_ (
);

AND2X2 _15732_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_4683_)
);

OR2X2 _15312_ (
    .A(_4265_),
    .B(_4268_),
    .Y(_4269_)
);

FILL FILL15200x301340 (
);

FILL FILL_0__10582_ (
);

BUFX2 BUFX2_insert40 (
    .A(_6289_),
    .Y(_6289__bF$buf4)
);

BUFX2 BUFX2_insert41 (
    .A(_6289_),
    .Y(_6289__bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .A(_6289_),
    .Y(_6289__bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .A(_6289_),
    .Y(_6289__bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .A(_6289_),
    .Y(_6289__bF$buf0)
);

BUFX2 BUFX2_insert45 (
    .A(_6310_),
    .Y(_6310__bF$buf4)
);

BUFX2 BUFX2_insert46 (
    .A(_6310_),
    .Y(_6310__bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .A(_6310_),
    .Y(_6310__bF$buf2)
);

FILL FILL319200x212420 (
);

BUFX2 BUFX2_insert48 (
    .A(_6310_),
    .Y(_6310__bF$buf1)
);

BUFX2 BUFX2_insert49 (
    .A(_6310_),
    .Y(_6310__bF$buf0)
);

FILL FILL_0__19280_ (
);

FILL FILL505400x227240 (
);

AND2X2 _16937_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_5869_)
);

AND2X2 _16517_ (
    .A(_4200__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_5455_)
);

FILL FILL_0__9381_ (
);

DFFSR _11652_ (
    .CLK(clk_bF$buf27),
    .D(_1587_[3]),
    .Q(\datapath_1.regfile_1.regOut[25] [3]),
    .R(rst_bF$buf28),
    .S(vdd)
);

FILL FILL_0__11367_ (
);

OR2X2 _11232_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_1433_)
);

OR2X2 _8859_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[4] [5]),
    .Y(_211_)
);

BUFX2 _8439_ (
    .A(_2_[15]),
    .Y(memoryWriteData[15])
);

FILL FILL372400x301340 (
);

FILL FILL180120x118560 (
);

AND2X2 _9800_ (
    .A(_698_),
    .B(_697_),
    .Y(_663_[17])
);

OR2X2 _12857_ (
    .A(_2421_),
    .B(_2419_),
    .Y(_2422_)
);

DFFSR _12437_ (
    .CLK(clk_bF$buf67),
    .D(_1983_[14]),
    .Q(\datapath_1.regfile_1.regOut[31] [14]),
    .R(rst_bF$buf60),
    .S(vdd)
);

AND2X2 _12017_ (
    .A(_1836_),
    .B(_1835_),
    .Y(_1785_[25])
);

FILL FILL145920x19760 (
);

FILL FILL_0__13513_ (
);

OR2X2 _16690_ (
    .A(_5624_),
    .B(_5625_),
    .Y(_5626_)
);

AND2X2 _16270_ (
    .A(_4208__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_5212_)
);

FILL FILL_1__9962_ (
);

FILL FILL_0__14718_ (
);

FILL FILL85120x123500 (
);

OR2X2 _17895_ (
    .A(_6799_),
    .B(_6812_),
    .Y(_6813_)
);

AND2X2 _17475_ (
    .A(_6399_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd1 [1])
);

OR2X2 _17055_ (
    .A(_5983_),
    .B(_5984_),
    .Y(_5985_)
);

DFFSR _12190_ (
    .CLK(clk_bF$buf69),
    .D(_1851_[25]),
    .Q(\datapath_1.regfile_1.regOut[29] [25]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL_0__18551_ (
);

FILL FILL_0__18131_ (
);

OR2X2 _9397_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .B(_530__bF$buf4),
    .Y(_490_)
);

FILL FILL_0__8652_ (
);

OR2X2 _10923_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_1267_)
);

FILL FILL_0__10218_ (
);

DFFSR _10503_ (
    .CLK(clk_bF$buf51),
    .D(_993_[15]),
    .Q(\datapath_1.regfile_1.regOut[16] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL20520x69160 (
);

FILL FILL237120x59280 (
);

XOR2X1 _13395_ (
    .A(_2393_),
    .B(_2931_),
    .Y(_2932_)
);

FILL FILL93480x237120 (
);

FILL FILL_0__19336_ (
);

OR2X2 _19201_ (
    .A(_8098_),
    .B(_8097_),
    .Y(_8099_)
);

FILL FILL_0__14891_ (
);

FILL FILL_0__9437_ (
);

AND2X2 _11708_ (
    .A(_1670_),
    .B(_1669_),
    .Y(_1653_[8])
);

FILL FILL351120x321100 (
);

FILL FILL_1__16263_ (
);

OR2X2 _15961_ (
    .A(_4907_),
    .B(_4892_),
    .Y(_4908_)
);

OR2X2 _15541_ (
    .A(_4493_),
    .B(_4494_),
    .Y(_4495_)
);

FILL FILL_0__15256_ (
);

FILL FILL64600x19760 (
);

AND2X2 _15121_ (
    .A(_4098_),
    .B(_4084_),
    .Y(_4099_)
);

FILL FILL90440x133380 (
);

FILL FILL_1__17468_ (
);

AND2X2 _16746_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_5681_)
);

AND2X2 _16326_ (
    .A(_4203__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_5267_)
);

OR2X2 _11881_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .B(_1784__bF$buf0),
    .Y(_1766_)
);

FILL FILL_0__9190_ (
);

OR2X2 _11461_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_1586__bF$buf3),
    .Y(_1546_)
);

FILL FILL_0__11176_ (
);

OR2X2 _11041_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .B(_1388__bF$buf4),
    .Y(_1326_)
);

FILL FILL_0__17402_ (
);

FILL FILL303240x242060 (
);

OR2X2 _8668_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_134__bF$buf2),
    .Y(_124_)
);

FILL FILL376960x217360 (
);

FILL FILL366320x177840 (
);

OR2X2 _12666_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(_2230_),
    .Y(_2231_)
);

OR2X2 _12246_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_1949_)
);

FILL FILL342760x83980 (
);

FILL FILL_0__18607_ (
);

FILL FILL_0__13742_ (
);

FILL FILL_0__13322_ (
);

FILL FILL106400x370500 (
);

FILL FILL19000x83980 (
);

FILL FILL_1__9771_ (
);

FILL FILL116280x316160 (
);

FILL FILL320720x118560 (
);

FILL FILL_1__15114_ (
);

FILL FILL_0__14947_ (
);

AND2X2 _14812_ (
    .A(_3907_),
    .B(_3906_),
    .Y(_3870_[18])
);

FILL FILL_0__14527_ (
);

FILL FILL_0__14107_ (
);

FILL FILL343520x202540 (
);

AND2X2 _17284_ (
    .A(_6203_),
    .B(_6209_),
    .Y(_6210_)
);

FILL FILL_0__18780_ (
);

FILL FILL_0__18360_ (
);

FILL FILL430160x113620 (
);

FILL FILL346560x83980 (
);

FILL FILL174040x103740 (
);

FILL FILL_0__8881_ (
);

FILL FILL_0__8461_ (
);

OR2X2 _10732_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_1190__bF$buf4),
    .Y(_1180_)
);

FILL FILL_0__10027_ (
);

OR2X2 _10312_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .B(_992__bF$buf3),
    .Y(_960_)
);

AND2X2 _18489_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_7398_)
);

AND2X2 _18069_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_6984_)
);

FILL FILL15960x247000 (
);

OR2X2 _19430_ (
    .A(gnd),
    .B(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_8322_)
);

OR2X2 _19010_ (
    .A(_7909_),
    .B(_7910_),
    .Y(_7911_)
);

FILL FILL_0__14280_ (
);

FILL FILL_0__9666_ (
);

DFFSR _11937_ (
    .CLK(clk_bF$buf70),
    .D(_1719_[30]),
    .Q(\datapath_1.regfile_1.regOut[27] [30]),
    .R(rst_bF$buf66),
    .S(vdd)
);

FILL FILL_0__9246_ (
);

OR2X2 _11517_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_1583_)
);

FILL FILL463600x29640 (
);

AND2X2 _15770_ (
    .A(_4236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_4720_)
);

FILL FILL_0__15485_ (
);

FILL FILL_0__15065_ (
);

OR2X2 _15350_ (
    .A(_4306_),
    .B(_4303_),
    .Y(_4307_)
);

FILL FILL12920x143260 (
);

FILL FILL_1__14805_ (
);

FILL FILL383800x44460 (
);

FILL FILL404320x316160 (
);

OR2X2 _16975_ (
    .A(_5905_),
    .B(_5904_),
    .Y(_5906_)
);

OR2X2 _16555_ (
    .A(_5492_),
    .B(_5491_),
    .Y(_5493_)
);

OR2X2 _16135_ (
    .A(_5077_),
    .B(_5078_),
    .Y(_5079_)
);

AND2X2 _11690_ (
    .A(_1658_),
    .B(_1657_),
    .Y(_1653_[2])
);

FILL FILL176320x44460 (
);

DFFSR _11270_ (
    .CLK(clk_bF$buf13),
    .D(_1389_[8]),
    .Q(\datapath_1.regfile_1.regOut[22] [8]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL360240x44460 (
);

FILL FILL_0__17631_ (
);

AND2X2 _8897_ (
    .A(_236_),
    .B(_235_),
    .Y(_201_[17])
);

AND2X2 _8477_ (
    .A(_16_),
    .B(_15_),
    .Y(_3_[6])
);

FILL FILL115520x167960 (
);

FILL FILL202920x172900 (
);

FILL FILL_1__10305_ (
);

FILL FILL380000x59280 (
);

FILL FILL_1__13197_ (
);

FILL FILL333640x291460 (
);

FILL FILL252320x227240 (
);

FILL FILL243200x83980 (
);

OR2X2 _12895_ (
    .A(_2458_),
    .B(_2459_),
    .Y(_2460_)
);

FILL FILL_1__19423_ (
);

OR2X2 _12475_ (
    .A(\aluControl_1.inst [4]),
    .B(_2067_),
    .Y(_2068_)
);

DFFSR _12055_ (
    .CLK(clk_bF$buf102),
    .D(_1785_[19]),
    .Q(\datapath_1.regfile_1.regOut[28] [19]),
    .R(rst_bF$buf41),
    .S(vdd)
);

FILL FILL304000x24700 (
);

OR2X2 _18701_ (
    .A(_7605_),
    .B(_7606_),
    .Y(_7607_)
);

FILL FILL_0__18416_ (
);

FILL FILL_0__13971_ (
);

FILL FILL387600x44460 (
);

FILL FILL_0__8937_ (
);

FILL FILL_1__9160_ (
);

FILL FILL_1__15763_ (
);

FILL FILL469680x24700 (
);

FILL FILL_0__14756_ (
);

FILL FILL146680x365560 (
);

DFFSR _14621_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[27]),
    .Q(\control_1.op [1]),
    .R(rst_bF$buf100),
    .S(vdd)
);

OR2X2 _14201_ (
    .A(\datapath_1.Data [19]),
    .B(_3605__bF$buf1),
    .Y(_3579_)
);

FILL FILL33440x167960 (
);

AND2X2 _17093_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_6022_)
);

FILL FILL387600x227240 (
);

FILL FILL489440x39520 (
);

FILL FILL56240x251940 (
);

AND2X2 _15826_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_4775_)
);

OR2X2 _15406_ (
    .A(_4360_),
    .B(_4361_),
    .Y(_4362_)
);

FILL FILL107920x182780 (
);

AND2X2 _10961_ (
    .A(_1292_),
    .B(_1291_),
    .Y(_1257_[17])
);

AND2X2 _10541_ (
    .A(_1072_),
    .B(_1071_),
    .Y(_1059_[6])
);

DFFSR _10121_ (
    .CLK(clk_bF$buf57),
    .D(_795_[20]),
    .Q(\datapath_1.regfile_1.regOut[13] [20]),
    .R(rst_bF$buf81),
    .S(vdd)
);

FILL FILL28880x286520 (
);

AND2X2 _18298_ (
    .A(_6236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_7210_)
);

FILL FILL_0__16902_ (
);

FILL FILL491720x148200 (
);

FILL FILL244720x242060 (
);

FILL FILL_0__19374_ (
);

FILL FILL_1__12468_ (
);

FILL FILL104880x227240 (
);

FILL FILL_0__9895_ (
);

OR2X2 _11746_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .B(_1718__bF$buf2),
    .Y(_1696_)
);

OR2X2 _11326_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .B(_1520__bF$buf3),
    .Y(_1476_)
);

FILL FILL130720x360620 (
);

FILL FILL_0__12822_ (
);

FILL FILL_0__12402_ (
);

FILL FILL199880x271700 (
);

FILL FILL127680x311220 (
);

FILL FILL_0__15294_ (
);

FILL FILL_1__8851_ (
);

FILL FILL191520x14820 (
);

FILL FILL_0__13607_ (
);

FILL FILL_1__17086_ (
);

FILL FILL248520x350740 (
);

OR2X2 _16784_ (
    .A(_5714_),
    .B(_5717_),
    .Y(_5718_)
);

AND2X2 _16364_ (
    .A(_4234__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_5305_)
);

FILL FILL354160x103740 (
);

FILL FILL434720x365560 (
);

FILL FILL_0__17860_ (
);

FILL FILL_0__17020_ (
);

BUFX2 BUFX2_insert480 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf0 )
);

BUFX2 BUFX2_insert481 (
    .A(_6250_),
    .Y(_6250__bF$buf4)
);

BUFX2 BUFX2_insert482 (
    .A(_6250_),
    .Y(_6250__bF$buf3)
);

BUFX2 BUFX2_insert483 (
    .A(_6250_),
    .Y(_6250__bF$buf2)
);

OR2X2 _17989_ (
    .A(_6904_),
    .B(_6905_),
    .Y(_6906_)
);

BUFX2 BUFX2_insert484 (
    .A(_6250_),
    .Y(_6250__bF$buf1)
);

OR2X2 _17569_ (
    .A(_6491_),
    .B(_6478_),
    .Y(_6492_)
);

BUFX2 BUFX2_insert485 (
    .A(_6250_),
    .Y(_6250__bF$buf0)
);

BUFX2 BUFX2_insert486 (
    .A(_3087_),
    .Y(_3087__bF$buf4)
);

OR2X2 _17149_ (
    .A(_6075_),
    .B(_6076_),
    .Y(_6077_)
);

BUFX2 BUFX2_insert487 (
    .A(_3087_),
    .Y(_3087__bF$buf3)
);

BUFX2 BUFX2_insert488 (
    .A(_3087_),
    .Y(_3087__bF$buf2)
);

BUFX2 BUFX2_insert489 (
    .A(_3087_),
    .Y(_3087__bF$buf1)
);

AND2X2 _12284_ (
    .A(_1974_),
    .B(_1973_),
    .Y(_1917_[28])
);

FILL FILL79800x118560 (
);

AND2X2 _18930_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_7832_)
);

FILL FILL_0__18225_ (
);

OR2X2 _18510_ (
    .A(_7415_),
    .B(_7418_),
    .Y(_7419_)
);

FILL FILL_0__13360_ (
);

FILL FILL_1__11739_ (
);

FILL FILL208240x34580 (
);

FILL FILL195320x14820 (
);

FILL FILL11400x59280 (
);

INVX2 _13489_ (
    .A(IorD_bF$buf3),
    .Y(_3079_)
);

NAND2X1 _13069_ (
    .A(_2524_),
    .B(_2624_),
    .Y(_2625_)
);

FILL FILL118560x69160 (
);

OR2X2 _14850_ (
    .A(\datapath_1.rd2 [31]),
    .B(_3935__bF$buf4),
    .Y(_3933_)
);

FILL FILL_0__14565_ (
);

FILL FILL_0__14145_ (
);

OR2X2 _14430_ (
    .A(memoryOutData[20]),
    .B(_3737__bF$buf2),
    .Y(_3713_)
);

AND2X2 _14010_ (
    .A(_3347__bF$buf0),
    .B(\datapath_1.PCJump [15]),
    .Y(_3428_)
);

FILL FILL328320x306280 (
);

FILL FILL_1__11492_ (
);

OR2X2 _15635_ (
    .A(_4585_),
    .B(_4586_),
    .Y(_4587_)
);

AND2X2 _15215_ (
    .A(_4172__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_4173_)
);

FILL FILL246240x212420 (
);

DFFSR _10770_ (
    .CLK(clk_bF$buf35),
    .D(_1125_[24]),
    .Q(\datapath_1.regfile_1.regOut[18] [24]),
    .R(rst_bF$buf67),
    .S(vdd)
);

FILL FILL_0__10065_ (
);

OR2X2 _10350_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_985_)
);

FILL FILL_0__16711_ (
);

FILL FILL384560x74100 (
);

AND2X2 _11975_ (
    .A(_1808_),
    .B(_1807_),
    .Y(_1785_[11])
);

FILL FILL_1__18923_ (
);

FILL FILL_0__9284_ (
);

AND2X2 _11555_ (
    .A(_1588_),
    .B(_1651_),
    .Y(_1587_[0])
);

DFFSR _11135_ (
    .CLK(clk_bF$buf111),
    .D(_1323_[2]),
    .Q(\datapath_1.regfile_1.regOut[21] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

FILL FILL_0__12631_ (
);

OR2X2 _9703_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .B(_662__bF$buf3),
    .Y(_654_)
);

FILL FILL202920x54340 (
);

FILL FILL_1__8660_ (
);

FILL FILL_1__14003_ (
);

FILL FILL468160x123500 (
);

FILL FILL_0__13836_ (
);

OR2X2 _13701_ (
    .A(_3180_),
    .B(_3179_),
    .Y(_3181_)
);

AND2X2 _16593_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_5530_)
);

AND2X2 _16173_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_5117_)
);

FILL FILL_1__15628_ (
);

OR2X2 _14906_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [7]),
    .Y(_3950_)
);

OR2X2 _17798_ (
    .A(_6686_),
    .B(_6717_),
    .Y(_6718_)
);

OR2X2 _17378_ (
    .A(_6303_),
    .B(_6301_),
    .Y(_6304_)
);

FILL FILL101080x167960 (
);

OR2X2 _12093_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_1867_)
);

FILL FILL198360x98800 (
);

FILL FILL382280x98800 (
);

FILL FILL_0__18874_ (
);

FILL FILL_0__18454_ (
);

FILL FILL_0__18034_ (
);

FILL FILL424840x108680 (
);

FILL FILL_0__8975_ (
);

AND2X2 _10826_ (
    .A(_1222_),
    .B(_1221_),
    .Y(_1191_[15])
);

AND2X2 _10406_ (
    .A(_1002_),
    .B(_1001_),
    .Y(_993_[4])
);

AND2X2 _13298_ (
    .A(_2839_),
    .B(_2838_),
    .Y(_2840_)
);

FILL FILL_0__11902_ (
);

FILL FILL_1__15381_ (
);

DFFSR _19524_ (
    .CLK(clk_bF$buf37),
    .D(_8320_[1]),
    .Q(\datapath_1.regfile_1.regOut[0] [1]),
    .R(rst_bF$buf87),
    .S(vdd)
);

AND2X2 _19104_ (
    .A(_6271__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_8003_)
);

FILL FILL_0__14374_ (
);

FILL FILL236360x167960 (
);

FILL FILL272840x340860 (
);

FILL FILL77520x59280 (
);

FILL FILL_1__16586_ (
);

OR2X2 _15864_ (
    .A(_4797_),
    .B(_4812_),
    .Y(_4813_)
);

FILL FILL_0__15579_ (
);

FILL FILL_0__15159_ (
);

AND2X2 _15444_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_4399_)
);

NOR2X1 _15024_ (
    .A(_4005_),
    .B(\datapath_1.a3 [2]),
    .Y(_4013_)
);

FILL FILL285000x74100 (
);

FILL FILL107160x158080 (
);

FILL FILL247000x19760 (
);

FILL FILL_0__16100_ (
);

FILL FILL189240x256880 (
);

FILL FILL67640x256880 (
);

OR2X2 _16649_ (
    .A(_5577_),
    .B(_5584_),
    .Y(_5585_)
);

AND2X2 _16229_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_5172_)
);

DFFSR _11784_ (
    .CLK(clk_bF$buf70),
    .D(_1653_[6]),
    .Q(\datapath_1.regfile_1.regOut[26] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

OR2X2 _11364_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_1501_)
);

FILL FILL_0__11079_ (
);

FILL FILL_0__17725_ (
);

FILL FILL_0__12860_ (
);

FILL FILL_0__12020_ (
);

AND2X2 _9932_ (
    .A(_766_),
    .B(_765_),
    .Y(_729_[18])
);

AND2X2 _9512_ (
    .A(_546_),
    .B(_545_),
    .Y(_531_[7])
);

OAI21X1 _12989_ (
    .A(_2500_),
    .B(_2322_),
    .C(_2383_),
    .Y(_2550_)
);

AND2X2 _12569_ (
    .A(_2089_),
    .B(_2108_),
    .Y(_2090_)
);

AND2X2 _12149_ (
    .A(_1904_),
    .B(_1903_),
    .Y(_1851_[26])
);

FILL FILL455240x0 (
);

FILL FILL_1__14652_ (
);

OR2X2 _13930_ (
    .A(_3359_),
    .B(_3358_),
    .Y(_3360_)
);

FILL FILL_0__13225_ (
);

OR2X2 _13510_ (
    .A(IorD_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [7]),
    .Y(_3028_)
);

BUFX2 BUFX2_insert1040 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf4 )
);

FILL FILL164920x128440 (
);

BUFX2 BUFX2_insert1041 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf3 )
);

BUFX2 BUFX2_insert1042 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf2 )
);

BUFX2 BUFX2_insert1043 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf1 )
);

BUFX2 BUFX2_insert1044 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf0 )
);

BUFX2 BUFX2_insert1045 (
    .A(_6328_),
    .Y(_6328__bF$buf4)
);

BUFX2 BUFX2_insert1046 (
    .A(_6328_),
    .Y(_6328__bF$buf3)
);

BUFX2 BUFX2_insert1047 (
    .A(_6328_),
    .Y(_6328__bF$buf2)
);

BUFX2 BUFX2_insert1048 (
    .A(_6328_),
    .Y(_6328__bF$buf1)
);

BUFX2 BUFX2_insert1049 (
    .A(_6328_),
    .Y(_6328__bF$buf0)
);

FILL FILL_1__10992_ (
);

FILL FILL145920x286520 (
);

OR2X2 _14715_ (
    .A(\datapath_1.rd1 [29]),
    .B(_3869__bF$buf3),
    .Y(_3863_)
);

BUFX2 BUFX2_insert860 (
    .A(_4230_),
    .Y(_4230__bF$buf2)
);

BUFX2 BUFX2_insert861 (
    .A(_4230_),
    .Y(_4230__bF$buf1)
);

BUFX2 BUFX2_insert862 (
    .A(_4230_),
    .Y(_4230__bF$buf0)
);

BUFX2 BUFX2_insert863 (
    .A(_266_),
    .Y(_266__bF$buf4)
);

BUFX2 BUFX2_insert864 (
    .A(_266_),
    .Y(_266__bF$buf3)
);

BUFX2 BUFX2_insert865 (
    .A(_266_),
    .Y(_266__bF$buf2)
);

BUFX2 BUFX2_insert866 (
    .A(_266_),
    .Y(_266__bF$buf1)
);

OR2X2 _17187_ (
    .A(_6113_),
    .B(_6114_),
    .Y(_6115_)
);

BUFX2 BUFX2_insert867 (
    .A(_266_),
    .Y(_266__bF$buf0)
);

BUFX2 BUFX2_insert868 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf4 )
);

BUFX2 BUFX2_insert869 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf3 )
);

FILL FILL_0__18683_ (
);

FILL FILL_0__8784_ (
);

DFFSR _10635_ (
    .CLK(clk_bF$buf110),
    .D(_1059_[18]),
    .Q(\datapath_1.regfile_1.regOut[17] [18]),
    .R(rst_bF$buf74),
    .S(vdd)
);

OR2X2 _10215_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_915_)
);

FILL FILL_0__11711_ (
);

FILL FILL_0__19468_ (
);

FILL FILL_0__19048_ (
);

OR2X2 _19333_ (
    .A(_8228_),
    .B(_8225_),
    .Y(_8229_)
);

FILL FILL_0__14183_ (
);

FILL FILL63840x286520 (
);

FILL FILL492480x113620 (
);

FILL FILL199880x39520 (
);

FILL FILL_1__13503_ (
);

FILL FILL505400x113620 (
);

FILL FILL401280x311220 (
);

FILL FILL_0__15388_ (
);

OR2X2 _15673_ (
    .A(_4624_),
    .B(_4593_),
    .Y(_4625_)
);

AND2X2 _15253_ (
    .A(_4210__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_4211_)
);

FILL FILL460560x9880 (
);

FILL FILL331360x316160 (
);

OR2X2 _16878_ (
    .A(_5810_),
    .B(_5809_),
    .Y(_5811_)
);

AND2X2 _16458_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_5397_)
);

OR2X2 _16038_ (
    .A(_4983_),
    .B(_4982_),
    .Y(_4984_)
);

OR2X2 _11593_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .B(_1652__bF$buf2),
    .Y(_1614_)
);

OR2X2 _11173_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .B(_1454__bF$buf3),
    .Y(_1394_)
);

FILL FILL142120x54340 (
);

FILL FILL_0__17954_ (
);

FILL FILL_0__17534_ (
);

FILL FILL_0__17114_ (
);

FILL FILL40280x217360 (
);

DFFSR _9741_ (
    .CLK(clk_bF$buf104),
    .D(_597_[27]),
    .Q(\datapath_1.regfile_1.regOut[10] [27]),
    .R(rst_bF$buf25),
    .S(vdd)
);

OR2X2 _9321_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_459_)
);

FILL FILL435480x330980 (
);

FILL FILL47120x93860 (
);

OR2X2 _12798_ (
    .A(_2362_),
    .B(_2350_),
    .Y(_2363_)
);

OR2X2 _12378_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_2017_)
);

FILL FILL_0__18739_ (
);

FILL FILL_0__18319_ (
);

OR2X2 _18604_ (
    .A(_7510_),
    .B(_7509_),
    .Y(_7511_)
);

FILL FILL297920x311220 (
);

FILL FILL_0__13874_ (
);

FILL FILL_0__13454_ (
);

FILL FILL_0__13034_ (
);

FILL FILL_1__9063_ (
);

FILL FILL83600x83980 (
);

FILL FILL278160x375440 (
);

AND2X2 _14944_ (
    .A(_3975_),
    .B(_3974_),
    .Y(_3936_[19])
);

FILL FILL_0__14659_ (
);

AND2X2 _14524_ (
    .A(_3755_),
    .B(_3754_),
    .Y(_3738_[8])
);

AND2X2 _14104_ (
    .A(_3352__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3509_)
);

FILL FILL183160x335920 (
);

FILL FILL67640x4940 (
);

FILL FILL_0__15600_ (
);

FILL FILL_0__18072_ (
);

FILL FILL_1__11166_ (
);

FILL FILL382280x296400 (
);

AND2X2 _15729_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_4680_)
);

AND2X2 _15309_ (
    .A(_4195__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_4266_)
);

FILL FILL_0__8593_ (
);

FILL FILL_0__10999_ (
);

OR2X2 _10864_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_1256__bF$buf3),
    .Y(_1248_)
);

FILL FILL_0__10159_ (
);

OR2X2 _10444_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .B(_1058__bF$buf2),
    .Y(_1028_)
);

FILL FILL505400x340860 (
);

OR2X2 _10024_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_860__bF$buf3),
    .Y(_808_)
);

FILL FILL_0__11940_ (
);

FILL FILL_0__11100_ (
);

AND2X2 _19142_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_8041_)
);

FILL FILL504640x59280 (
);

FILL FILL491720x39520 (
);

FILL FILL_0__9798_ (
);

DFFSR _11649_ (
    .CLK(clk_bF$buf99),
    .D(_1587_[0]),
    .Q(\datapath_1.regfile_1.regOut[25] [0]),
    .R(rst_bF$buf19),
    .S(vdd)
);

OR2X2 _11229_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_1431_)
);

FILL FILL_1__13732_ (
);

FILL FILL308560x276640 (
);

FILL FILL53960x163020 (
);

FILL FILL_0__12725_ (
);

FILL FILL129960x34580 (
);

AND2X2 _15482_ (
    .A(_4436_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.rd2 [3])
);

AND2X2 _15062_ (
    .A(_4048_),
    .B(_4050_),
    .Y(_4051_)
);

FILL FILL_1__8754_ (
);

FILL FILL_1__14937_ (
);

FILL FILL376960x103740 (
);

OR2X2 _16687_ (
    .A(_5619_),
    .B(_5622_),
    .Y(_5623_)
);

AND2X2 _16267_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_5209_)
);

FILL FILL_1__18350_ (
);

FILL FILL406600x153140 (
);

FILL FILL_1__9119_ (
);

FILL FILL_0__17343_ (
);

FILL FILL_1__10437_ (
);

OR2X2 _9970_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_794__bF$buf4),
    .Y(_792_)
);

OR2X2 _9550_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .B(_596__bF$buf1),
    .Y(_572_)
);

OR2X2 _9130_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .B(_398__bF$buf0),
    .Y(_352_)
);

FILL FILL442320x232180 (
);

FILL FILL393680x340860 (
);

FILL FILL_1__19555_ (
);

DFFSR _12187_ (
    .CLK(clk_bF$buf26),
    .D(_1851_[22]),
    .Q(\datapath_1.regfile_1.regOut[29] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL_0__18968_ (
);

FILL FILL_0__18548_ (
);

AND2X2 _18833_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_7737_)
);

FILL FILL_0_BUFX2_insert500 (
);

FILL FILL_0_BUFX2_insert501 (
);

OR2X2 _18413_ (
    .A(_7315_),
    .B(_7322_),
    .Y(_7323_)
);

FILL FILL_0_BUFX2_insert502 (
);

FILL FILL_0_BUFX2_insert503 (
);

FILL FILL342000x326040 (
);

FILL FILL_0__13683_ (
);

FILL FILL_0_BUFX2_insert505 (
);

FILL FILL_0__13263_ (
);

FILL FILL_0_BUFX2_insert507 (
);

FILL FILL228000x350740 (
);

FILL FILL_0_BUFX2_insert509 (
);

FILL FILL444600x9880 (
);

FILL FILL_1__15055_ (
);

FILL FILL68400x143260 (
);

FILL FILL_1__10190_ (
);

FILL FILL_0__14888_ (
);

DFFSR _14753_ (
    .CLK(clk_bF$buf40),
    .D(_3804_[30]),
    .Q(\datapath_1.a [30]),
    .R(rst_bF$buf63),
    .S(vdd)
);

FILL FILL_0__14048_ (
);

OR2X2 _14333_ (
    .A(vdd),
    .B(ALUOut[31]),
    .Y(_3668_)
);

FILL FILL440800x266760 (
);

FILL FILL210520x34580 (
);

FILL FILL463600x9880 (
);

FILL FILL437760x217360 (
);

FILL FILL427120x177840 (
);

OR2X2 _15958_ (
    .A(_4903_),
    .B(_4904_),
    .Y(_4905_)
);

OR2X2 _15538_ (
    .A(_4491_),
    .B(_4490_),
    .Y(_4492_)
);

AND2X2 _15118_ (
    .A(_4096_),
    .B(_4095_),
    .Y(_4097_)
);

FILL FILL108680x14820 (
);

AND2X2 _10673_ (
    .A(_1140_),
    .B(_1139_),
    .Y(_1125_[7])
);

DFFSR _10253_ (
    .CLK(clk_bF$buf101),
    .D(_861_[23]),
    .Q(\datapath_1.regfile_1.regOut[14] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL_0__16614_ (
);

AND2X2 _19371_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_8266_)
);

FILL FILL_0__19086_ (
);

DFFSR _8821_ (
    .CLK(clk_bF$buf107),
    .D(_135_[10]),
    .Q(\datapath_1.regfile_1.regOut[3] [10]),
    .R(rst_bF$buf95),
    .S(vdd)
);

BUFX2 _8401_ (
    .A(_1_[9]),
    .Y(memoryAddress[9])
);

OR2X2 _11878_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .B(_1784__bF$buf0),
    .Y(_1764_)
);

FILL FILL_0__9187_ (
);

OR2X2 _11458_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .B(_1586__bF$buf2),
    .Y(_1544_)
);

OR2X2 _11038_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_1388__bF$buf1),
    .Y(_1324_)
);

FILL FILL_1__13121_ (
);

FILL FILL_0__17819_ (
);

FILL FILL_0__12954_ (
);

FILL FILL_0__12534_ (
);

FILL FILL164920x19760 (
);

AND2X2 _15291_ (
    .A(_4203__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_4248_)
);

DFFSR _9606_ (
    .CLK(clk_bF$buf106),
    .D(_531_[21]),
    .Q(\datapath_1.regfile_1.regOut[9] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

FILL FILL_0__13739_ (
);

FILL FILL_0__13319_ (
);

OR2X2 _13604_ (
    .A(_3097_),
    .B(_3094_),
    .Y(\datapath_1.mux_pcsrc.dout [1])
);

AND2X2 _16496_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_5435_)
);

OR2X2 _16076_ (
    .A(_5020_),
    .B(_5019_),
    .Y(_5021_)
);

FILL FILL47120x163020 (
);

FILL FILL_0__17992_ (
);

FILL FILL_0__17572_ (
);

FILL FILL_0__17152_ (
);

FILL FILL182400x118560 (
);

AND2X2 _14809_ (
    .A(_3905_),
    .B(_3904_),
    .Y(_3870_[17])
);

FILL FILL168720x19760 (
);

FILL FILL_1__19364_ (
);

FILL FILL_0__10600_ (
);

OR2X2 _18642_ (
    .A(_7533_),
    .B(_7548_),
    .Y(_7549_)
);

AND2X2 _18222_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_7135_)
);

FILL FILL442320x370500 (
);

FILL FILL_0__13072_ (
);

FILL FILL319960x271700 (
);

FILL FILL_0__8878_ (
);

OR2X2 _10729_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .B(_1190__bF$buf4),
    .Y(_1178_)
);

OR2X2 _10309_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_992__bF$buf4),
    .Y(_958_)
);

FILL FILL283480x311220 (
);

FILL FILL9120x123500 (
);

INVX2 _19427_ (
    .A(gnd),
    .Y(_8385_)
);

FILL FILL87400x123500 (
);

OR2X2 _19007_ (
    .A(_7904_),
    .B(_7907_),
    .Y(_7908_)
);

FILL FILL_0__14697_ (
);

DFFSR _14982_ (
    .CLK(clk_bF$buf62),
    .D(_3936_[1]),
    .Q(\datapath_1.mux_iord.din0 [1]),
    .R(rst_bF$buf18),
    .S(vdd)
);

OR2X2 _14562_ (
    .A(memoryOutData[21]),
    .B(_3803__bF$buf4),
    .Y(_3781_)
);

FILL FILL_0__14277_ (
);

OR2X2 _14142_ (
    .A(ALUOut[0]),
    .B(MemToReg_bF$buf3),
    .Y(_3604_)
);

FILL FILL_1__16069_ (
);

OR2X2 _15767_ (
    .A(_4716_),
    .B(_4713_),
    .Y(_4717_)
);

AND2X2 _15347_ (
    .A(_4135__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_4304_)
);

FILL FILL_0__10197_ (
);

OR2X2 _10482_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_1053_)
);

OR2X2 _10062_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_833_)
);

FILL FILL_1__17010_ (
);

FILL FILL_0__16843_ (
);

FILL FILL_0__16423_ (
);

FILL FILL_0__16003_ (
);

FILL FILL129200x256880 (
);

OR2X2 _19180_ (
    .A(_8070_),
    .B(_8077_),
    .Y(_8078_)
);

FILL FILL298680x167960 (
);

AND2X2 _8630_ (
    .A(_98_),
    .B(_97_),
    .Y(_69_[14])
);

FILL FILL30400x247000 (
);

FILL FILL353400x321100 (
);

AND2X2 _11687_ (
    .A(_1656_),
    .B(_1655_),
    .Y(_1653_[1])
);

FILL FILL_1__18215_ (
);

DFFSR _11267_ (
    .CLK(clk_bF$buf29),
    .D(_1389_[5]),
    .Q(\datapath_1.regfile_1.regOut[22] [5]),
    .R(rst_bF$buf48),
    .S(vdd)
);

AND2X2 _17913_ (
    .A(_6262__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_6831_)
);

FILL FILL_0__17208_ (
);

FILL FILL_0__12343_ (
);

FILL FILL408880x118560 (
);

OR2X2 _9835_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .B(_728__bF$buf2),
    .Y(_722_)
);

OR2X2 _9415_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .B(_530__bF$buf0),
    .Y(_502_)
);

FILL FILL_1__8792_ (
);

FILL FILL92720x133380 (
);

FILL FILL_1__14555_ (
);

FILL FILL484120x306280 (
);

FILL FILL_0__13548_ (
);

AND2X2 _13833_ (
    .A(_3288_),
    .B(_3287_),
    .Y(\datapath_1.alu_1.ALUInA [5])
);

FILL FILL_0__13128_ (
);

AND2X2 _13413_ (
    .A(_2948_),
    .B(_2937_),
    .Y(_2949_)
);

FILL FILL298680x44460 (
);

FILL FILL451440x167960 (
);

FILL FILL387600x340860 (
);

FILL FILL279680x113620 (
);

DFFSR _14618_ (
    .CLK(clk_bF$buf65),
    .D(_3738_[24]),
    .Q(\datapath_1.PCJump [26]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _18871_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_7774_)
);

FILL FILL_0__18586_ (
);

FILL FILL_0__18166_ (
);

AND2X2 _18451_ (
    .A(_6300__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_7360_)
);

OR2X2 _18031_ (
    .A(_6945_),
    .B(_6946_),
    .Y(_6947_)
);

FILL FILL118560x316160 (
);

AND2X2 _10958_ (
    .A(_1290_),
    .B(_1289_),
    .Y(_1257_[16])
);

AND2X2 _10538_ (
    .A(_1070_),
    .B(_1069_),
    .Y(_1059_[5])
);

DFFSR _10118_ (
    .CLK(clk_bF$buf64),
    .D(_795_[17]),
    .Q(\datapath_1.regfile_1.regOut[13] [17]),
    .R(rst_bF$buf10),
    .S(vdd)
);

FILL FILL_1__12621_ (
);

FILL FILL104880x340860 (
);

FILL FILL_0__11614_ (
);

FILL FILL22800x128440 (
);

OR2X2 _19236_ (
    .A(_8131_),
    .B(_8132_),
    .Y(_8133_)
);

AND2X2 _14791_ (
    .A(_3893_),
    .B(_3892_),
    .Y(_3870_[11])
);

AND2X2 _14371_ (
    .A(_3673_),
    .B(_3736_),
    .Y(_3672_[0])
);

FILL FILL345040x108680 (
);

FILL FILL432440x113620 (
);

FILL FILL156560x4940 (
);

FILL FILL176320x103740 (
);

FILL FILL275120x29640 (
);

FILL FILL165680x49400 (
);

FILL FILL_0__12819_ (
);

FILL FILL413440x271700 (
);

AND2X2 _15996_ (
    .A(_4177__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_4942_)
);

OR2X2 _15576_ (
    .A(_4521_),
    .B(_4528_),
    .Y(_4529_)
);

NOR2X1 _15156_ (
    .A(_4119_),
    .B(_4042_),
    .Y(\datapath_1.regfile_1.regEn [26])
);

OR2X2 _10291_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_992__bF$buf1),
    .Y(_946_)
);

FILL FILL_0__16652_ (
);

FILL FILL174800x271700 (
);

FILL FILL_1__18864_ (
);

OR2X2 _11496_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[24] [24]),
    .Y(_1569_)
);

FILL FILL_1__18444_ (
);

OR2X2 _11076_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_1349_)
);

FILL FILL_0__17437_ (
);

OR2X2 _17722_ (
    .A(_6642_),
    .B(_6641_),
    .Y(_6643_)
);

AND2X2 _17302_ (
    .A(_6226_),
    .B(_6227_),
    .Y(_6228_)
);

FILL FILL_0__17017_ (
);

FILL FILL226480x345800 (
);

FILL FILL_0__12992_ (
);

FILL FILL_0__12572_ (
);

FILL FILL_0__12152_ (
);

AND2X2 _9644_ (
    .A(_614_),
    .B(_613_),
    .Y(_597_[8])
);

DFFSR _9224_ (
    .CLK(clk_bF$buf54),
    .D(_333_[26]),
    .Q(\datapath_1.regfile_1.regOut[6] [26]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL437000x93860 (
);

FILL FILL_1__19229_ (
);

FILL FILL406600x316160 (
);

AND2X2 _18927_ (
    .A(_6317__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_7829_)
);

AND2X2 _18507_ (
    .A(_6238__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_7416_)
);

FILL FILL_0__13777_ (
);

OR2X2 _13642_ (
    .A(_3128_),
    .B(_3129_),
    .Y(_3130_)
);

NOR2X1 _13222_ (
    .A(_2503_),
    .B(_2214_),
    .Y(_2769_)
);

FILL FILL318440x281580 (
);

FILL FILL237120x217360 (
);

FILL FILL_0__17190_ (
);

FILL FILL_1__15569_ (
);

FILL FILL_1__15149_ (
);

FILL FILL335920x291460 (
);

FILL FILL350360x163020 (
);

FILL FILL254600x227240 (
);

OR2X2 _14847_ (
    .A(\datapath_1.rd2 [30]),
    .B(_3935__bF$buf1),
    .Y(_3931_)
);

OR2X2 _14427_ (
    .A(memoryOutData[19]),
    .B(_3737__bF$buf3),
    .Y(_3711_)
);

OR2X2 _14007_ (
    .A(_3425_),
    .B(_3424_),
    .Y(_3426_)
);

FILL FILL_1__16510_ (
);

FILL FILL_0_CLKBUF1_insert110 (
);

FILL FILL_0_CLKBUF1_insert111 (
);

FILL FILL_0_CLKBUF1_insert113 (
);

FILL FILL_0_CLKBUF1_insert115 (
);

FILL FILL_0_CLKBUF1_insert117 (
);

FILL FILL_0_CLKBUF1_insert119 (
);

FILL FILL277400x311220 (
);

AND2X2 _18680_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_7586_)
);

FILL FILL_0__18395_ (
);

AND2X2 _18260_ (
    .A(_6312__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_7172_)
);

FILL FILL5320x9880 (
);

FILL FILL_0__8496_ (
);

DFFSR _10767_ (
    .CLK(clk_bF$buf47),
    .D(_1125_[21]),
    .Q(\datapath_1.regfile_1.regOut[18] [21]),
    .R(rst_bF$buf103),
    .S(vdd)
);

OR2X2 _10347_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_983_)
);

FILL FILL_1__12850_ (
);

FILL FILL_1__12010_ (
);

FILL FILL_0__16708_ (
);

FILL FILL_0__11843_ (
);

FILL FILL_0__11423_ (
);

FILL FILL35720x167960 (
);

AND2X2 _19465_ (
    .A(_8345_),
    .B(_8344_),
    .Y(_8320_[12])
);

FILL FILL304000x98800 (
);

OR2X2 _19045_ (
    .A(_7943_),
    .B(_7944_),
    .Y(_7945_)
);

FILL FILL341240x74100 (
);

OR2X2 _14180_ (
    .A(\datapath_1.Data [12]),
    .B(_3605__bF$buf2),
    .Y(_3565_)
);

FILL FILL459040x128440 (
);

FILL FILL273600x49400 (
);

AND2X2 _8915_ (
    .A(_248_),
    .B(_247_),
    .Y(_201_[23])
);

FILL FILL384560x182780 (
);

FILL FILL6080x192660 (
);

FILL FILL_1_BUFX2_insert431 (
);

NOR2X1 _12913_ (
    .A(_2321_),
    .B(_2325_),
    .Y(_2478_)
);

FILL FILL_0__12208_ (
);

FILL FILL_1_BUFX2_insert433 (
);

FILL FILL_1_BUFX2_insert435 (
);

FILL FILL12160x232180 (
);

OR2X2 _15385_ (
    .A(_4340_),
    .B(_4325_),
    .Y(_4341_)
);

FILL FILL499320x222300 (
);

FILL FILL_0__16461_ (
);

FILL FILL_0__16041_ (
);

BUFX2 BUFX2_insert100 (
    .A(_1850_),
    .Y(_1850__bF$buf4)
);

BUFX2 BUFX2_insert101 (
    .A(_1850_),
    .Y(_1850__bF$buf3)
);

FILL FILL129960x311220 (
);

BUFX2 BUFX2_insert102 (
    .A(_1850_),
    .Y(_1850__bF$buf2)
);

BUFX2 BUFX2_insert103 (
    .A(_1850_),
    .Y(_1850__bF$buf1)
);

FILL FILL_0__17666_ (
);

AND2X2 _17951_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_6868_)
);

BUFX2 BUFX2_insert104 (
    .A(_1850_),
    .Y(_1850__bF$buf0)
);

BUFX2 BUFX2_insert105 (
    .A(IorD),
    .Y(IorD_bF$buf4)
);

OR2X2 _17531_ (
    .A(_6453_),
    .B(_6454_),
    .Y(_6455_)
);

BUFX2 BUFX2_insert106 (
    .A(IorD),
    .Y(IorD_bF$buf3)
);

OR2X2 _17111_ (
    .A(_6036_),
    .B(_6039_),
    .Y(_6040_)
);

BUFX2 BUFX2_insert107 (
    .A(IorD),
    .Y(IorD_bF$buf2)
);

BUFX2 BUFX2_insert108 (
    .A(IorD),
    .Y(IorD_bF$buf1)
);

FILL FILL_0__12381_ (
);

BUFX2 BUFX2_insert109 (
    .A(IorD),
    .Y(IorD_bF$buf0)
);

FILL FILL196840x9880 (
);

DFFSR _9873_ (
    .CLK(clk_bF$buf54),
    .D(_663_[30]),
    .Q(\datapath_1.regfile_1.regOut[11] [30]),
    .R(rst_bF$buf48),
    .S(vdd)
);

OR2X2 _9453_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_527_)
);

OR2X2 _9033_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_307_)
);

FILL FILL_1__11701_ (
);

FILL FILL326800x59280 (
);

FILL FILL_1__14173_ (
);

AND2X2 _18736_ (
    .A(_6250__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_7641_)
);

OR2X2 _18316_ (
    .A(_7220_),
    .B(_7227_),
    .Y(_7228_)
);

OR2X2 _13871_ (
    .A(\datapath_1.a [18]),
    .B(_3342__bF$buf4),
    .Y(_3314_)
);

FILL FILL_0__13166_ (
);

AND2X2 _13451_ (
    .A(_2664_),
    .B(_2695_),
    .Y(_2984_)
);

OR2X2 _13031_ (
    .A(_2157__bF$buf2),
    .B(_2588_),
    .Y(_2589_)
);

FILL FILL408880x39520 (
);

FILL FILL_1__9195_ (
);

FILL FILL50920x360620 (
);

FILL FILL_0__9913_ (
);

FILL FILL_1__15798_ (
);

FILL FILL47880x311220 (
);

FILL FILL474240x321100 (
);

AND2X2 _14656_ (
    .A(_3823_),
    .B(_3822_),
    .Y(_3804_[9])
);

OR2X2 _14236_ (
    .A(MemToReg_bF$buf1),
    .B(ALUOut[31]),
    .Y(_3602_)
);

FILL FILL_0__15732_ (
);

FILL FILL_0__15312_ (
);

FILL FILL390640x350740 (
);

FILL FILL_1__11298_ (
);

OR2X2 _10996_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_1322__bF$buf3),
    .Y(_1316_)
);

OR2X2 _10576_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .B(_1124__bF$buf2),
    .Y(_1096_)
);

OR2X2 _10156_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_926__bF$buf3),
    .Y(_876_)
);

FILL FILL196080x74100 (
);

FILL FILL_0__16937_ (
);

FILL FILL_0__16517_ (
);

AND2X2 _16802_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_5736_)
);

FILL FILL_0__11232_ (
);

OR2X2 _19274_ (
    .A(_8169_),
    .B(_8170_),
    .Y(_8171_)
);

OR2X2 _8724_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_141_)
);

FILL FILL_1__18729_ (
);

FILL FILL_1__18309_ (
);

FILL FILL417240x217360 (
);

FILL FILL_0__12857_ (
);

OR2X2 _12722_ (
    .A(_2286_),
    .B(_2259_),
    .Y(_2287_)
);

DFFSR _12302_ (
    .CLK(clk_bF$buf67),
    .D(_1917_[8]),
    .Q(\datapath_1.regfile_1.regOut[30] [8]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_0__12017_ (
);

FILL FILL261440x207480 (
);

FILL FILL299440x0 (
);

AND2X2 _15194_ (
    .A(_4151__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_4152_)
);

AND2X2 _9929_ (
    .A(_764_),
    .B(_763_),
    .Y(_729_[17])
);

AND2X2 _9509_ (
    .A(_544_),
    .B(_543_),
    .Y(_531_[6])
);

FILL FILL_1__8886_ (
);

FILL FILL229520x370500 (
);

FILL FILL_0__16690_ (
);

FILL FILL_0__16270_ (
);

OR2X2 _13927_ (
    .A(_3355_),
    .B(_3356_),
    .Y(_3357_)
);

OR2X2 _13507_ (
    .A(IorD_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [6]),
    .Y(_3026_)
);

FILL FILL85880x345800 (
);

OR2X2 _16399_ (
    .A(_5337_),
    .B(_5338_),
    .Y(_5339_)
);

FILL FILL_1__18482_ (
);

AND2X2 _17760_ (
    .A(_6247__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_6680_)
);

FILL FILL_0__17055_ (
);

OR2X2 _17340_ (
    .A(_6265_),
    .B(_6263_),
    .Y(_6266_)
);

FILL FILL_1__10569_ (
);

FILL FILL396720x207480 (
);

FILL FILL263720x296400 (
);

OR2X2 _9682_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .B(_662__bF$buf0),
    .Y(_640_)
);

FILL FILL269040x370500 (
);

OR2X2 _9262_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .B(_464__bF$buf2),
    .Y(_420_)
);

FILL FILL_1_CLKBUF1_insert141 (
);

FILL FILL202160x54340 (
);

FILL FILL_0__10923_ (
);

FILL FILL96520x217360 (
);

OR2X2 _18965_ (
    .A(_7863_),
    .B(_7866_),
    .Y(_7867_)
);

OR2X2 _18545_ (
    .A(_7452_),
    .B(_7439_),
    .Y(_7453_)
);

AND2X2 _18125_ (
    .A(_7039_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.rd1 [11])
);

FILL FILL_0__13395_ (
);

OR2X2 _13680_ (
    .A(_3162_),
    .B(_3161_),
    .Y(_3163_)
);

XOR2X1 _13260_ (
    .A(_2221_),
    .B(_2804_),
    .Y(_2805_)
);

FILL FILL_0__19201_ (
);

FILL FILL_1__12715_ (
);

FILL FILL_0__11708_ (
);

FILL FILL_0__9302_ (
);

FILL FILL481840x286520 (
);

FILL FILL_1__15187_ (
);

INVX2 _14885_ (
    .A(PCEn_bF$buf1),
    .Y(_4001_)
);

DFFSR _14465_ (
    .CLK(clk_bF$buf65),
    .D(_3672_[0]),
    .Q(\datapath_1.Data [0]),
    .R(rst_bF$buf26),
    .S(vdd)
);

AND2X2 _14045_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3458_)
);

FILL FILL103360x167960 (
);

FILL FILL_0__15961_ (
);

FILL FILL_0__15541_ (
);

FILL FILL_0__15121_ (
);

DFFSR _10385_ (
    .CLK(clk_bF$buf86),
    .D(_927_[26]),
    .Q(\datapath_1.regfile_1.regOut[15] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

FILL FILL_1__17333_ (
);

FILL FILL380000x108680 (
);

OR2X2 _16611_ (
    .A(_5547_),
    .B(_5546_),
    .Y(_5548_)
);

FILL FILL_0__11461_ (
);

FILL FILL361000x266760 (
);

AND2X2 _19083_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_7983_)
);

FILL FILL238640x167960 (
);

DFFSR _8953_ (
    .CLK(clk_bF$buf85),
    .D(_201_[13]),
    .Q(\datapath_1.regfile_1.regOut[4] [13]),
    .R(rst_bF$buf60),
    .S(vdd)
);

OR2X2 _8533_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .B(_68__bF$buf4),
    .Y(_54_)
);

FILL FILL71440x316160 (
);

FILL FILL_1__18958_ (
);

FILL FILL_1__13673_ (
);

OR2X2 _17816_ (
    .A(_6727_),
    .B(_6734_),
    .Y(_6735_)
);

FILL FILL_1_BUFX2_insert811 (
);

XOR2X1 _12951_ (
    .A(_2356_),
    .B(_2513_),
    .Y(_2514_)
);

FILL FILL_0__12666_ (
);

FILL FILL_1_BUFX2_insert813 (
);

AND2X2 _12531_ (
    .A(\control_1.op [0]),
    .B(\control_1.op [1]),
    .Y(_2121_)
);

OR2X2 _12111_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_1879_)
);

FILL FILL_1_BUFX2_insert815 (
);

FILL FILL109440x158080 (
);

DFFSR _9738_ (
    .CLK(clk_bF$buf97),
    .D(_597_[24]),
    .Q(\datapath_1.regfile_1.regOut[10] [24]),
    .R(rst_bF$buf84),
    .S(vdd)
);

FILL FILL462080x138320 (
);

OR2X2 _9318_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_457_)
);

FILL FILL291840x256880 (
);

FILL FILL69920x256880 (
);

FILL FILL_1__14038_ (
);

OR2X2 _13736_ (
    .A(_3210_),
    .B(_3209_),
    .Y(_3211_)
);

AND2X2 _13316_ (
    .A(_2392_),
    .B(_2393_),
    .Y(_2857_)
);

FILL FILL_0__14812_ (
);

FILL FILL101080x350740 (
);

FILL FILL_0__17284_ (
);

AND2X2 _9491_ (
    .A(_532_),
    .B(_595_),
    .Y(_531_[0])
);

DFFSR _9071_ (
    .CLK(clk_bF$buf112),
    .D(_267_[2]),
    .Q(\datapath_1.regfile_1.regOut[5] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

FILL FILL_0__10732_ (
);

FILL FILL_0__10312_ (
);

OR2X2 _18774_ (
    .A(_7645_),
    .B(_7678_),
    .Y(_7679_)
);

FILL FILL_0__18489_ (
);

FILL FILL13680x182780 (
);

OR2X2 _18354_ (
    .A(_7263_),
    .B(_7264_),
    .Y(_7265_)
);

FILL FILL_0__19430_ (
);

FILL FILL_1__17809_ (
);

FILL FILL183920x83980 (
);

FILL FILL_0__9531_ (
);

FILL FILL_0__9111_ (
);

DFFSR _11802_ (
    .CLK(clk_bF$buf35),
    .D(_1653_[24]),
    .Q(\datapath_1.regfile_1.regOut[26] [24]),
    .R(rst_bF$buf6),
    .S(vdd)
);

OR2X2 _19559_ (
    .A(_8389_),
    .B(_8387_),
    .Y(PCEn)
);

AND2X2 _19139_ (
    .A(_6326__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_8038_)
);

FILL FILL253840x360620 (
);

OR2X2 _14694_ (
    .A(\datapath_1.rd1 [22]),
    .B(_3869__bF$buf2),
    .Y(_3849_)
);

OR2X2 _14274_ (
    .A(\datapath_1.ALUResult [11]),
    .B(_3671__bF$buf2),
    .Y(_3629_)
);

FILL FILL_0__15770_ (
);

AND2X2 _15899_ (
    .A(_4151__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_4847_)
);

OR2X2 _15479_ (
    .A(_4433_),
    .B(_4426_),
    .Y(_4434_)
);

OR2X2 _15059_ (
    .A(\datapath_1.a3 [4]),
    .B(_4021_),
    .Y(_4048_)
);

FILL FILL_1__17982_ (
);

FILL FILL_1__17562_ (
);

OR2X2 _10194_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_901_)
);

FILL FILL221920x98800 (
);

FILL FILL_0__16555_ (
);

OR2X2 _16840_ (
    .A(_5769_),
    .B(_5772_),
    .Y(_5773_)
);

FILL FILL_0__16135_ (
);

AND2X2 _16420_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_5360_)
);

OR2X2 _16000_ (
    .A(_4944_),
    .B(_4945_),
    .Y(_4946_)
);

FILL FILL_0__11690_ (
);

AND2X2 _8762_ (
    .A(_166_),
    .B(_165_),
    .Y(_135_[15])
);

FILL FILL114000x177840 (
);

DFFSR _11399_ (
    .CLK(clk_bF$buf63),
    .D(_1455_[8]),
    .Q(\datapath_1.regfile_1.regOut[23] [8]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL_1__13062_ (
);

OR2X2 _17625_ (
    .A(_6546_),
    .B(_6545_),
    .Y(_6547_)
);

FILL FILL403560x311220 (
);

OR2X2 _17205_ (
    .A(_6132_),
    .B(_6131_),
    .Y(_6133_)
);

FILL FILL_0__12895_ (
);

OR2X2 _12760_ (
    .A(_2324_),
    .B(_2323_),
    .Y(_2325_)
);

FILL FILL_0__12475_ (
);

FILL FILL418760x0 (
);

OR2X2 _12340_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .B(_2048__bF$buf2),
    .Y(_1992_)
);

FILL FILL_0__18701_ (
);

OR2X2 _9967_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .B(_794__bF$buf0),
    .Y(_790_)
);

FILL FILL333640x316160 (
);

OR2X2 _9547_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_596__bF$buf0),
    .Y(_570_)
);

OR2X2 _9127_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_398__bF$buf2),
    .Y(_350_)
);

FILL FILL234080x212420 (
);

FILL FILL_1__14687_ (
);

FILL FILL_0_BUFX2_insert470 (
);

FILL FILL_0_BUFX2_insert472 (
);

FILL FILL_0_BUFX2_insert474 (
);

OR2X2 _13965_ (
    .A(_3389_),
    .B(_3388_),
    .Y(_3390_)
);

FILL FILL245480x281580 (
);

AND2X2 _13545_ (
    .A(_3051_),
    .B(_3050_),
    .Y(_1_[18])
);

FILL FILL_0_BUFX2_insert475 (
);

OR2X2 _13125_ (
    .A(_2677_),
    .B(_2449_),
    .Y(_2678_)
);

FILL FILL_0_BUFX2_insert476 (
);

FILL FILL_0_BUFX2_insert477 (
);

FILL FILL_0_BUFX2_insert478 (
);

FILL FILL251560x222300 (
);

FILL FILL_0__14201_ (
);

FILL FILL42560x217360 (
);

FILL FILL_0__17093_ (
);

FILL FILL65360x301340 (
);

FILL FILL300200x301340 (
);

FILL FILL_0__15826_ (
);

FILL FILL_0__15406_ (
);

FILL FILL_0__10961_ (
);

FILL FILL_0__10541_ (
);

OR2X2 _18583_ (
    .A(_7488_),
    .B(_7489_),
    .Y(_7490_)
);

AND2X2 _18163_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_7077_)
);

FILL FILL103360x237120 (
);

FILL FILL_0__11746_ (
);

OR2X2 _11611_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .B(_1652__bF$buf0),
    .Y(_1626_)
);

AND2X2 _19368_ (
    .A(_6321__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_8263_)
);

FILL FILL185440x335920 (
);

AND2X2 _14083_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3491_)
);

FILL FILL367080x286520 (
);

DFFSR _8818_ (
    .CLK(clk_bF$buf66),
    .D(_135_[7]),
    .Q(\datapath_1.regfile_1.regOut[3] [7]),
    .R(rst_bF$buf80),
    .S(vdd)
);

FILL FILL120840x247000 (
);

FILL FILL148960x34580 (
);

FILL FILL_1__13538_ (
);

OAI21X1 _12816_ (
    .A(_2158_),
    .B(_2376__bF$buf3),
    .C(_2380_),
    .Y(_2381_)
);

OR2X2 _15288_ (
    .A(_4245_),
    .B(_4221_),
    .Y(_4246_)
);

FILL FILL_0__16784_ (
);

FILL FILL_1__9501_ (
);

OR2X2 _8991_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_279_)
);

DFFSR _8571_ (
    .CLK(clk_bF$buf37),
    .D(_3_[18]),
    .Q(\datapath_1.regfile_1.regOut[1] [18]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL325280x148200 (
);

FILL FILL_1__13291_ (
);

FILL FILL416480x350740 (
);

FILL FILL361760x321100 (
);

FILL FILL_0__17569_ (
);

AND2X2 _17854_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_6773_)
);

OR2X2 _17434_ (
    .A(_6357_),
    .B(_6358_),
    .Y(_6359_)
);

FILL FILL_0__17149_ (
);

OR2X2 _17014_ (
    .A(_5941_),
    .B(_5944_),
    .Y(_5945_)
);

FILL FILL_0__12284_ (
);

FILL FILL_0__18930_ (
);

FILL FILL291840x326040 (
);

AND2X2 _9776_ (
    .A(_682_),
    .B(_681_),
    .Y(_663_[9])
);

DFFSR _9356_ (
    .CLK(clk_bF$buf0),
    .D(_399_[29]),
    .Q(\datapath_1.regfile_1.regOut[7] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

FILL FILL_0__8611_ (
);

FILL FILL158840x187720 (
);

OR2X2 _18639_ (
    .A(_7544_),
    .B(_7545_),
    .Y(_7546_)
);

OR2X2 _18219_ (
    .A(_7131_),
    .B(_7118_),
    .Y(_7132_)
);

AND2X2 _13774_ (
    .A(_3084__bF$buf2),
    .B(\datapath_1.PCJump [26]),
    .Y(_3243_)
);

FILL FILL_0__13489_ (
);

INVX1 _13354_ (
    .A(_2406_),
    .Y(_2893_)
);

FILL FILL_0__14850_ (
);

FILL FILL_0__14010_ (
);

FILL FILL_0__9816_ (
);

FILL FILL395960x340860 (
);

FILL FILL78280x340860 (
);

OR2X2 _14979_ (
    .A(\datapath_1.mux_pcsrc.dout [31]),
    .B(_4001__bF$buf4),
    .Y(_3999_)
);

OR2X2 _14559_ (
    .A(memoryOutData[20]),
    .B(_3803__bF$buf4),
    .Y(_3779_)
);

AND2X2 _14139_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3539_)
);

FILL FILL304760x217360 (
);

FILL FILL_0__15635_ (
);

AND2X2 _15920_ (
    .A(_4236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_4868_)
);

OR2X2 _15500_ (
    .A(_4453_),
    .B(_4452_),
    .Y(_4454_)
);

FILL FILL_0__10350_ (
);

OR2X2 _18392_ (
    .A(_7298_),
    .B(_7301_),
    .Y(_7302_)
);

FILL FILL256120x291460 (
);

DFFSR _10899_ (
    .CLK(clk_bF$buf6),
    .D(_1191_[24]),
    .Q(\datapath_1.regfile_1.regOut[19] [24]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL_1__17847_ (
);

FILL FILL_1__17427_ (
);

OR2X2 _10479_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_1051_)
);

OR2X2 _10059_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_831_)
);

FILL FILL_1__12142_ (
);

OR2X2 _16705_ (
    .A(_5639_),
    .B(_5636_),
    .Y(_5640_)
);

FILL FILL107160x79040 (
);

FILL FILL_0__11975_ (
);

AND2X2 _11840_ (
    .A(_1738_),
    .B(_1737_),
    .Y(_1719_[9])
);

DFFSR _11420_ (
    .CLK(clk_bF$buf88),
    .D(_1455_[29]),
    .Q(\datapath_1.regfile_1.regOut[23] [29]),
    .R(rst_bF$buf112),
    .S(vdd)
);

AND2X2 _11000_ (
    .A(_1318_),
    .B(_1317_),
    .Y(_1257_[30])
);

AND2X2 _19177_ (
    .A(_6293__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_8075_)
);

AND2X2 _8627_ (
    .A(_96_),
    .B(_95_),
    .Y(_69_[13])
);

FILL FILL429400x177840 (
);

FILL FILL325280x375440 (
);

FILL FILL408120x44460 (
);

XNOR2X1 _12625_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2190_)
);

OR2X2 _12205_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .B(_1982__bF$buf4),
    .Y(_1922_)
);

NAND3X1 _15097_ (
    .A(_4018_),
    .B(\datapath_1.a3 [3]),
    .C(_4019_),
    .Y(_4080_)
);

FILL FILL_0__13701_ (
);

FILL FILL_0__16173_ (
);

FILL FILL_1__9310_ (
);

FILL FILL_0__14906_ (
);

FILL FILL130720x182780 (
);

FILL FILL127680x133380 (
);

FILL FILL108680x88920 (
);

FILL FILL_0__17798_ (
);

AND2X2 _17663_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_6585_)
);

FILL FILL_0__17378_ (
);

AND2X2 _17243_ (
    .A(_4241__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_6170_)
);

FILL FILL_0__12093_ (
);

DFFSR _9585_ (
    .CLK(clk_bF$buf99),
    .D(_531_[0]),
    .Q(\datapath_1.regfile_1.regOut[9] [0]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9165_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_375_)
);

FILL FILL_1__11833_ (
);

FILL FILL_0__8420_ (
);

FILL FILL504640x182780 (
);

FILL FILL_0__10406_ (
);

OR2X2 _18868_ (
    .A(_7763_),
    .B(_7770_),
    .Y(_7771_)
);

FILL FILL_0_BUFX2_insert850 (
);

OR2X2 _18448_ (
    .A(_7325_),
    .B(_7357_),
    .Y(_7358_)
);

FILL FILL_0_BUFX2_insert852 (
);

OR2X2 _18028_ (
    .A(_6942_),
    .B(_6943_),
    .Y(_6944_)
);

FILL FILL_0_BUFX2_insert854 (
);

FILL FILL_0__13298_ (
);

OR2X2 _13583_ (
    .A(ALUOut[31]),
    .B(_3079__bF$buf3),
    .Y(_3077_)
);

FILL FILL_0_BUFX2_insert855 (
);

AND2X2 _13163_ (
    .A(_2713_),
    .B(_2701_),
    .Y(_2714_)
);

FILL FILL_0_BUFX2_insert856 (
);

FILL FILL_0_BUFX2_insert857 (
);

FILL FILL_0_BUFX2_insert858 (
);

FILL FILL446120x202540 (
);

FILL FILL_0__9625_ (
);

AND2X2 _14788_ (
    .A(_3891_),
    .B(_3890_),
    .Y(_3870_[10])
);

OR2X2 _14368_ (
    .A(\datapath_1.Data [0]),
    .B(vdd),
    .Y(_3736_)
);

FILL FILL_1__16451_ (
);

FILL FILL_1__16031_ (
);

FILL FILL262960x227240 (
);

FILL FILL_0__15024_ (
);

BUFX2 BUFX2_insert10 (
    .A(_3344_),
    .Y(_3344__bF$buf4)
);

BUFX2 BUFX2_insert11 (
    .A(_3344_),
    .Y(_3344__bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .A(_3344_),
    .Y(_3344__bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .A(_3344_),
    .Y(_3344__bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .A(_3344_),
    .Y(_3344__bF$buf0)
);

BUFX2 BUFX2_insert15 (
    .A(_4167_),
    .Y(_4167__bF$buf4)
);

BUFX2 BUFX2_insert16 (
    .A(_4167_),
    .Y(_4167__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .A(_4167_),
    .Y(_4167__bF$buf2)
);

FILL FILL198360x306280 (
);

BUFX2 BUFX2_insert18 (
    .A(_4167_),
    .Y(_4167__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .A(_4167_),
    .Y(_4167__bF$buf0)
);

FILL FILL57000x375440 (
);

FILL FILL295640x34580 (
);

OR2X2 _10288_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_992__bF$buf1),
    .Y(_944_)
);

FILL FILL_1__12791_ (
);

FILL FILL_0__16649_ (
);

OR2X2 _16934_ (
    .A(_5864_),
    .B(_5865_),
    .Y(_5866_)
);

AND2X2 _16514_ (
    .A(_4189__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_5452_)
);

FILL FILL_0__16229_ (
);

FILL FILL_0__11364_ (
);

OR2X2 _8856_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_209_)
);

BUFX2 _8436_ (
    .A(_2_[12]),
    .Y(memoryWriteData[12])
);

FILL FILL_1__13156_ (
);

OR2X2 _17719_ (
    .A(_6638_),
    .B(_6639_),
    .Y(_6640_)
);

FILL FILL66880x251940 (
);

FILL FILL_0__12989_ (
);

NAND3X1 _12854_ (
    .A(_2416_),
    .B(_2417_),
    .C(_2418_),
    .Y(_2419_)
);

DFFSR _12434_ (
    .CLK(clk_bF$buf79),
    .D(_1983_[11]),
    .Q(\datapath_1.regfile_1.regOut[31] [11]),
    .R(rst_bF$buf12),
    .S(vdd)
);

AND2X2 _12014_ (
    .A(_1834_),
    .B(_1833_),
    .Y(_1785_[24])
);

FILL FILL333640x49400 (
);

FILL FILL_0__13930_ (
);

FILL FILL227240x192660 (
);

FILL FILL237120x330980 (
);

FILL FILL319200x148200 (
);

FILL FILL216600x88920 (
);

OR2X2 _13639_ (
    .A(_3127_),
    .B(_3124_),
    .Y(\datapath_1.mux_pcsrc.dout [6])
);

XOR2X1 _13219_ (
    .A(_2214_),
    .B(_2765_),
    .Y(_2766_)
);

FILL FILL230280x64220 (
);

OR2X2 _17892_ (
    .A(_6808_),
    .B(_6809_),
    .Y(_6810_)
);

OR2X2 _17472_ (
    .A(_6381_),
    .B(_6396_),
    .Y(_6397_)
);

OR2X2 _17052_ (
    .A(_5981_),
    .B(_5980_),
    .Y(_5982_)
);

FILL FILL280440x281580 (
);

FILL FILL_1__16927_ (
);

OR2X2 _9394_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .B(_530__bF$buf3),
    .Y(_488_)
);

FILL FILL180120x375440 (
);

FILL FILL_1__11642_ (
);

FILL FILL_1__19399_ (
);

FILL FILL177080x326040 (
);

OR2X2 _10920_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_1265_)
);

DFFSR _10500_ (
    .CLK(clk_bF$buf60),
    .D(_993_[12]),
    .Q(\datapath_1.regfile_1.regOut[16] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

AND2X2 _18677_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_7583_)
);

AND2X2 _18257_ (
    .A(_6264__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_7169_)
);

NAND2X1 _13392_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2929_)
);

FILL FILL_0__19333_ (
);

FILL FILL453720x167960 (
);

FILL FILL_0__9434_ (
);

FILL FILL_0__9014_ (
);

AND2X2 _11705_ (
    .A(_1668_),
    .B(_1667_),
    .Y(_1653_[7])
);

FILL FILL346560x4940 (
);

DFFSR _14597_ (
    .CLK(clk_bF$buf23),
    .D(_3738_[3]),
    .Q(\aluControl_1.inst [3]),
    .R(rst_bF$buf22),
    .S(vdd)
);

OR2X2 _14177_ (
    .A(\datapath_1.Data [11]),
    .B(_3605__bF$buf3),
    .Y(_3563_)
);

FILL FILL_1__16680_ (
);

FILL FILL155800x153140 (
);

FILL FILL_0__15673_ (
);

FILL FILL_0__15253_ (
);

FILL FILL376200x345800 (
);

FILL FILL298680x350740 (
);

FILL FILL251560x88920 (
);

AND2X2 _10097_ (
    .A(_856_),
    .B(_855_),
    .Y(_795_[30])
);

FILL FILL_0__16878_ (
);

OR2X2 _16743_ (
    .A(_5674_),
    .B(_5677_),
    .Y(_5678_)
);

FILL FILL_0__16038_ (
);

AND2X2 _16323_ (
    .A(_4236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_5264_)
);

FILL FILL_0__11593_ (
);

FILL FILL_0__11173_ (
);

OR2X2 _8665_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .B(_134__bF$buf2),
    .Y(_122_)
);

FILL FILL178600x103740 (
);

AND2X2 _17948_ (
    .A(_6250__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_6865_)
);

FILL FILL73720x153140 (
);

OR2X2 _17528_ (
    .A(_6451_),
    .B(_6448_),
    .Y(_6452_)
);

AND2X2 _17108_ (
    .A(_4181__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_6037_)
);

FILL FILL_0__12798_ (
);

FILL FILL41800x365560 (
);

OR2X2 _12663_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(_2227_),
    .Y(_2228_)
);

OR2X2 _12243_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_1947_)
);

FILL FILL237880x59280 (
);

OR2X2 _13868_ (
    .A(\datapath_1.a [17]),
    .B(_3342__bF$buf0),
    .Y(_3312_)
);

AND2X2 _13448_ (
    .A(_2977_),
    .B(_2980_),
    .Y(_2981_)
);

AND2X2 _13028_ (
    .A(_2575_),
    .B(_2586_),
    .Y(_2587_)
);

FILL FILL117040x163020 (
);

FILL FILL193800x187720 (
);

AND2X2 _17281_ (
    .A(_6206__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_6207_)
);

FILL FILL_1__16316_ (
);

FILL FILL_1__11451_ (
);

FILL FILL_0__10864_ (
);

FILL FILL_0__10444_ (
);

AND2X2 _18486_ (
    .A(_6328__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_7395_)
);

AND2X2 _18066_ (
    .A(_6328__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_6981_)
);

FILL FILL_0__19142_ (
);

FILL FILL_1__12656_ (
);

FILL FILL352640x163020 (
);

FILL FILL_0__9243_ (
);

DFFSR _11934_ (
    .CLK(clk_bF$buf59),
    .D(_1719_[27]),
    .Q(\datapath_1.regfile_1.regOut[27] [27]),
    .R(rst_bF$buf92),
    .S(vdd)
);

OR2X2 _11514_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_1581_)
);

AND2X2 _12719_ (
    .A(_2282_),
    .B(_2283_),
    .Y(_2284_)
);

FILL FILL_1_BUFX2_insert76 (
);

FILL FILL_1_BUFX2_insert78 (
);

FILL FILL19760x83980 (
);

FILL FILL_0__16687_ (
);

OR2X2 _16972_ (
    .A(_5902_),
    .B(_5901_),
    .Y(_5903_)
);

OR2X2 _16552_ (
    .A(_5489_),
    .B(_5482_),
    .Y(_5490_)
);

FILL FILL_0__16267_ (
);

FILL FILL364040x74100 (
);

OR2X2 _16132_ (
    .A(_5074_),
    .B(_5075_),
    .Y(_5076_)
);

FILL FILL_1__9404_ (
);

AND2X2 _8894_ (
    .A(_234_),
    .B(_233_),
    .Y(_201_[16])
);

FILL FILL75240x123500 (
);

AND2X2 _8474_ (
    .A(_14_),
    .B(_13_),
    .Y(_3_[5])
);

FILL FILL_1__10722_ (
);

FILL FILL_1__18899_ (
);

AND2X2 _17757_ (
    .A(_6321__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_6677_)
);

FILL FILL14440x232180 (
);

FILL FILL401280x133380 (
);

AND2X2 _17337_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_6263_)
);

NAND2X1 _12892_ (
    .A(_2280_),
    .B(_2288_),
    .Y(_2457_)
);

FILL FILL366320x9880 (
);

AND2X2 _12472_ (
    .A(_2064_),
    .B(_2061_),
    .Y(_2065_)
);

DFFSR _12052_ (
    .CLK(clk_bF$buf78),
    .D(_1785_[16]),
    .Q(\datapath_1.regfile_1.regOut[28] [16]),
    .R(rst_bF$buf110),
    .S(vdd)
);

FILL FILL345800x59280 (
);

FILL FILL_0__18833_ (
);

FILL FILL_0__18413_ (
);

FILL FILL231800x326040 (
);

OR2X2 _9679_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_662__bF$buf2),
    .Y(_638_)
);

OR2X2 _9259_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .B(_464__bF$buf4),
    .Y(_418_)
);

FILL FILL_0__8514_ (
);

FILL FILL390640x197600 (
);

OR2X2 _13677_ (
    .A(_3158_),
    .B(_3159_),
    .Y(_3160_)
);

FILL FILL349600x4940 (
);

AND2X2 _13257_ (
    .A(_2801_),
    .B(_2433_),
    .Y(_2802_)
);

FILL FILL_1_BUFX2_insert1166 (
);

FILL FILL_1_BUFX2_insert1168 (
);

AND2X2 _17090_ (
    .A(_4208__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_6019_)
);

FILL FILL33440x44460 (
);

FILL FILL271320x326040 (
);

FILL FILL368600x4940 (
);

FILL FILL_1__16965_ (
);

FILL FILL_1__16545_ (
);

FILL FILL349600x59280 (
);

FILL FILL436240x0 (
);

FILL FILL297920x133380 (
);

FILL FILL_0__15538_ (
);

OR2X2 _15823_ (
    .A(_4771_),
    .B(_4770_),
    .Y(_4772_)
);

FILL FILL_0__15118_ (
);

OR2X2 _15403_ (
    .A(_4357_),
    .B(_4358_),
    .Y(_4359_)
);

FILL FILL_0__10673_ (
);

FILL FILL422560x251940 (
);

AND2X2 _18295_ (
    .A(_6326__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_7207_)
);

FILL FILL_0__19371_ (
);

OR2X2 _16608_ (
    .A(_5541_),
    .B(_5544_),
    .Y(_5545_)
);

FILL FILL_0__11878_ (
);

FILL FILL_0__11458_ (
);

OR2X2 _11743_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .B(_1718__bF$buf3),
    .Y(_1694_)
);

FILL FILL_0__9052_ (
);

OR2X2 _11323_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .B(_1520__bF$buf3),
    .Y(_1474_)
);

FILL FILL_0__11038_ (
);

FILL FILL52440x266760 (
);

FILL FILL380760x59280 (
);

FILL FILL_0__15291_ (
);

FILL FILL243960x83980 (
);

INVX1 _12948_ (
    .A(_2511_),
    .Y(\datapath_1.ALUResult [30])
);

AND2X2 _12528_ (
    .A(_2096_),
    .B(_2117_),
    .Y(_2118_)
);

OR2X2 _12108_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_1877_)
);

FILL FILL_1_BUFX2_insert786 (
);

FILL FILL_1_BUFX2_insert788 (
);

FILL FILL_0__13604_ (
);

FILL FILL_0__16496_ (
);

AND2X2 _16781_ (
    .A(_4195__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_5715_)
);

FILL FILL_0__16076_ (
);

AND2X2 _16361_ (
    .A(_4189__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_5302_)
);

FILL FILL_1__10531_ (
);

FILL FILL_0__14809_ (
);

FILL FILL_1__18288_ (
);

BUFX2 BUFX2_insert450 (
    .A(_1256_),
    .Y(_1256__bF$buf0)
);

BUFX2 BUFX2_insert451 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf4 )
);

BUFX2 BUFX2_insert452 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf3 )
);

BUFX2 BUFX2_insert453 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf2 )
);

BUFX2 BUFX2_insert454 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf1 )
);

OR2X2 _17986_ (
    .A(_6901_),
    .B(_6902_),
    .Y(_6903_)
);

OR2X2 _17566_ (
    .A(_6488_),
    .B(_6487_),
    .Y(_6489_)
);

BUFX2 BUFX2_insert455 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf0 )
);

BUFX2 BUFX2_insert456 (
    .A(_4225_),
    .Y(_4225__bF$buf4)
);

AND2X2 _17146_ (
    .A(_6074_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd2 [29])
);

BUFX2 BUFX2_insert457 (
    .A(_4225_),
    .Y(_4225__bF$buf3)
);

BUFX2 BUFX2_insert458 (
    .A(_4225_),
    .Y(_4225__bF$buf2)
);

BUFX2 BUFX2_insert459 (
    .A(_4225_),
    .Y(_4225__bF$buf1)
);

AND2X2 _12281_ (
    .A(_1972_),
    .B(_1971_),
    .Y(_1917_[27])
);

FILL FILL_0__18642_ (
);

FILL FILL244720x365560 (
);

OR2X2 _9488_ (
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .Y(_595_)
);

AND2X2 _9068_ (
    .A(_330_),
    .B(_329_),
    .Y(_267_[31])
);

FILL FILL181640x113620 (
);

FILL FILL_0__8743_ (
);

FILL FILL_0__10729_ (
);

FILL FILL_0__10309_ (
);

OR2X2 _13486_ (
    .A(\datapath_1.PCJump_17_bF$buf2 ),
    .B(_3005_),
    .Y(_3014_)
);

AND2X2 _13066_ (
    .A(_2622_),
    .B(_2607_),
    .Y(_2623_)
);

FILL FILL504640x296400 (
);

FILL FILL468920x202540 (
);

FILL FILL_0__19427_ (
);

FILL FILL_0__19007_ (
);

FILL FILL_0__14562_ (
);

FILL FILL_0__14142_ (
);

FILL FILL_0__9948_ (
);

FILL FILL_0__9528_ (
);

FILL FILL299440x103740 (
);

FILL FILL449160x266760 (
);

FILL FILL157320x29640 (
);

FILL FILL_0__15767_ (
);

FILL FILL_0__15347_ (
);

OR2X2 _15632_ (
    .A(_4580_),
    .B(_4583_),
    .Y(_4584_)
);

INVX1 _15212_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_4170_)
);

FILL FILL_0__10482_ (
);

FILL FILL_0__10062_ (
);

FILL FILL367080x172900 (
);

FILL FILL_0__19180_ (
);

FILL FILL80560x271700 (
);

FILL FILL459800x54340 (
);

FILL FILL306280x281580 (
);

FILL FILL297160x177840 (
);

AND2X2 _16837_ (
    .A(_4172__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_5770_)
);

FILL FILL155800x316160 (
);

AND2X2 _16417_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_5357_)
);

FILL FILL312360x222300 (
);

FILL FILL_0__9281_ (
);

AND2X2 _11972_ (
    .A(_1806_),
    .B(_1805_),
    .Y(_1785_[10])
);

FILL FILL105640x167960 (
);

OR2X2 _11552_ (
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .Y(_1651_)
);

AND2X2 _11132_ (
    .A(_1386_),
    .B(_1385_),
    .Y(_1323_[31])
);

FILL FILL281200x59280 (
);

FILL FILL_0__17913_ (
);

AND2X2 _8759_ (
    .A(_164_),
    .B(_163_),
    .Y(_135_[14])
);

FILL FILL242440x227240 (
);

FILL FILL456000x69160 (
);

OR2X2 _9700_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .B(_662__bF$buf1),
    .Y(_652_)
);

FILL FILL_1__13479_ (
);

NAND2X1 _12757_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2322_)
);

OR2X2 _12337_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .B(_2048__bF$buf2),
    .Y(_1990_)
);

FILL FILL_1__14840_ (
);

FILL FILL56240x306280 (
);

FILL FILL_0__13413_ (
);

AND2X2 _16590_ (
    .A(_4197__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_5527_)
);

AND2X2 _16170_ (
    .A(_4135__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_5114_)
);

FILL FILL_1__9442_ (
);

FILL FILL386080x158080 (
);

OR2X2 _14903_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [6]),
    .Y(_3948_)
);

FILL FILL291080x118560 (
);

OR2X2 _17795_ (
    .A(_6711_),
    .B(_6714_),
    .Y(_6715_)
);

AND2X2 _17375_ (
    .A(_6300__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_6301_)
);

OR2X2 _12090_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_1865_)
);

FILL FILL_0__18451_ (
);

FILL FILL_0__18031_ (
);

OR2X2 _9297_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_443_)
);

FILL FILL_0__8972_ (
);

FILL FILL_0__8552_ (
);

AND2X2 _10823_ (
    .A(_1220_),
    .B(_1219_),
    .Y(_1191_[14])
);

FILL FILL_0__10538_ (
);

AND2X2 _10403_ (
    .A(_1000_),
    .B(_999_),
    .Y(_993_[3])
);

OR2X2 _13295_ (
    .A(_2157__bF$buf3),
    .B(_2836_),
    .Y(_2837_)
);

FILL FILL103360x350740 (
);

FILL FILL287280x54340 (
);

OR2X2 _19521_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8383_)
);

FILL FILL_0__19236_ (
);

AND2X2 _19101_ (
    .A(_6206__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_8000_)
);

FILL FILL_0__14791_ (
);

FILL FILL_0__14371_ (
);

FILL FILL387600x0 (
);

FILL FILL_0__9757_ (
);

OR2X2 _11608_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .B(_1652__bF$buf2),
    .Y(_1624_)
);

FILL FILL_0__15996_ (
);

OR2X2 _15861_ (
    .A(_4809_),
    .B(_4808_),
    .Y(_4810_)
);

FILL FILL_0__15156_ (
);

AND2X2 _15441_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_4396_)
);

NAND3X1 _15021_ (
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .C(\datapath_1.a3 [4]),
    .Y(_4010_)
);

FILL FILL_0__10291_ (
);

FILL FILL342000x286520 (
);

FILL FILL21280x350740 (
);

FILL FILL267520x24700 (
);

FILL FILL_1__17368_ (
);

FILL FILL183160x227240 (
);

AND2X2 _16646_ (
    .A(_4130__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_5582_)
);

AND2X2 _16226_ (
    .A(_4195__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_5169_)
);

DFFSR _11781_ (
    .CLK(clk_bF$buf46),
    .D(_1653_[3]),
    .Q(\datapath_1.regfile_1.regOut[26] [3]),
    .R(rst_bF$buf97),
    .S(vdd)
);

FILL FILL_0__11496_ (
);

OR2X2 _11361_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_1499_)
);

FILL FILL_0__17302_ (
);

OR2X2 _8988_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_277_)
);

DFFSR _8568_ (
    .CLK(clk_bF$buf90),
    .D(_3_[15]),
    .Q(\datapath_1.regfile_1.regOut[1] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL505400x232180 (
);

FILL FILL272840x276640 (
);

INVX1 _12986_ (
    .A(_2387__bF$buf1),
    .Y(_2547_)
);

AND2X2 _12566_ (
    .A(_2085_),
    .B(_2086_),
    .Y(_2087_)
);

AND2X2 _12146_ (
    .A(_1902_),
    .B(_1901_),
    .Y(_1851_[25])
);

FILL FILL_0__18927_ (
);

FILL FILL_0__18507_ (
);

FILL FILL_0__13642_ (
);

FILL FILL_0__8608_ (
);

FILL FILL_1__9251_ (
);

BUFX2 BUFX2_insert1010 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf4 )
);

BUFX2 BUFX2_insert1011 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf3 )
);

BUFX2 BUFX2_insert1012 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf2 )
);

BUFX2 BUFX2_insert1013 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf1 )
);

BUFX2 BUFX2_insert1014 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf0 )
);

BUFX2 BUFX2_insert1015 (
    .A(_3935_),
    .Y(_3935__bF$buf4)
);

BUFX2 BUFX2_insert1016 (
    .A(_3935_),
    .Y(_3935__bF$buf3)
);

BUFX2 BUFX2_insert1017 (
    .A(_3935_),
    .Y(_3935__bF$buf2)
);

FILL FILL_1__15434_ (
);

BUFX2 BUFX2_insert1018 (
    .A(_3935_),
    .Y(_3935__bF$buf1)
);

FILL FILL_1__15014_ (
);

BUFX2 BUFX2_insert1019 (
    .A(_3935_),
    .Y(_3935__bF$buf0)
);

FILL FILL405840x311220 (
);

FILL FILL_0__14847_ (
);

OR2X2 _14712_ (
    .A(\datapath_1.rd1 [28]),
    .B(_3869__bF$buf2),
    .Y(_3861_)
);

FILL FILL_0__14427_ (
);

FILL FILL_0__14007_ (
);

BUFX2 BUFX2_insert830 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf2 )
);

BUFX2 BUFX2_insert831 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf1 )
);

BUFX2 BUFX2_insert832 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf0 )
);

BUFX2 BUFX2_insert833 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf4)
);

BUFX2 BUFX2_insert834 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf3)
);

BUFX2 BUFX2_insert835 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf2)
);

BUFX2 BUFX2_insert836 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf1)
);

OR2X2 _17184_ (
    .A(_6108_),
    .B(_6111_),
    .Y(_6112_)
);

BUFX2 BUFX2_insert837 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf0)
);

BUFX2 BUFX2_insert838 (
    .A(_134_),
    .Y(_134__bF$buf4)
);

BUFX2 BUFX2_insert839 (
    .A(_134_),
    .Y(_134__bF$buf3)
);

FILL FILL_0__18680_ (
);

FILL FILL_0__18260_ (
);

FILL FILL_1__11774_ (
);

AND2X2 _15917_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_4865_)
);

FILL FILL217360x370500 (
);

FILL FILL247760x281580 (
);

FILL FILL247760x19760 (
);

DFFSR _10632_ (
    .CLK(clk_bF$buf112),
    .D(_1059_[15]),
    .Q(\datapath_1.regfile_1.regOut[17] [15]),
    .R(rst_bF$buf3),
    .S(vdd)
);

OR2X2 _10212_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_913_)
);

FILL FILL253840x222300 (
);

AND2X2 _18389_ (
    .A(_6323__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_7299_)
);

AND2X2 _19330_ (
    .A(_6289__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_8226_)
);

FILL FILL_0__14180_ (
);

FILL FILL_0__9566_ (
);

AND2X2 _11837_ (
    .A(_1736_),
    .B(_1735_),
    .Y(_1719_[8])
);

FILL FILL_0__9146_ (
);

DFFSR _11417_ (
    .CLK(clk_bF$buf30),
    .D(_1455_[26]),
    .Q(\datapath_1.regfile_1.regOut[23] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL_1__13920_ (
);

FILL FILL_0__12913_ (
);

FILL FILL_0__15385_ (
);

OR2X2 _15670_ (
    .A(_4621_),
    .B(_4618_),
    .Y(_4622_)
);

AND2X2 _15250_ (
    .A(_4207_),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .Y(_4208_)
);

FILL FILL461320x172900 (
);

FILL FILL209760x0 (
);

FILL FILL_1__8522_ (
);

FILL FILL469680x192660 (
);

FILL FILL97280x163020 (
);

FILL FILL105640x237120 (
);

OR2X2 _16875_ (
    .A(_5806_),
    .B(_5807_),
    .Y(_5808_)
);

OR2X2 _16455_ (
    .A(_5393_),
    .B(_5392_),
    .Y(_5394_)
);

OR2X2 _16035_ (
    .A(_4980_),
    .B(_4979_),
    .Y(_4981_)
);

FILL FILL211280x311220 (
);

OR2X2 _11590_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .B(_1652__bF$buf0),
    .Y(_1612_)
);

OR2X2 _11170_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .B(_1454__bF$buf2),
    .Y(_1392_)
);

FILL FILL369360x286520 (
);

FILL FILL_0__17951_ (
);

FILL FILL_0__17531_ (
);

OR2X2 _8797_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .B(_200__bF$buf3),
    .Y(_190_)
);

FILL FILL15200x123500 (
);

FILL FILL386840x296400 (
);

FILL FILL107920x54340 (
);

FILL FILL_1__13097_ (
);

INVX1 _12795_ (
    .A(_2359_),
    .Y(_2360_)
);

OR2X2 _12375_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_2015_)
);

FILL FILL_0__18316_ (
);

OR2X2 _18601_ (
    .A(_7503_),
    .B(_7507_),
    .Y(_7508_)
);

FILL FILL_0__13871_ (
);

FILL FILL_0__13031_ (
);

FILL FILL_0__8417_ (
);

FILL FILL480320x158080 (
);

FILL FILL503120x29640 (
);

FILL FILL285000x118560 (
);

FILL FILL372400x123500 (
);

FILL FILL_1__15663_ (
);

FILL FILL_0__14656_ (
);

AND2X2 _14941_ (
    .A(_3973_),
    .B(_3972_),
    .Y(_3936_[18])
);

FILL FILL_0__14236_ (
);

AND2X2 _14521_ (
    .A(_3753_),
    .B(_3752_),
    .Y(_3738_[7])
);

AND2X2 _14101_ (
    .A(_3347__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3506_)
);

FILL FILL262960x340860 (
);

FILL FILL_1__11583_ (
);

OR2X2 _15726_ (
    .A(_4675_),
    .B(_4676_),
    .Y(_4677_)
);

FILL FILL63080x237120 (
);

AND2X2 _15306_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_4263_)
);

FILL FILL386080x311220 (
);

FILL FILL_0__10996_ (
);

FILL FILL_0__10576_ (
);

OR2X2 _10861_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .B(_1256__bF$buf0),
    .Y(_1246_)
);

OR2X2 _10441_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .B(_1058__bF$buf2),
    .Y(_1026_)
);

OR2X2 _10021_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_860__bF$buf3),
    .Y(_806_)
);

AND2X2 _18198_ (
    .A(_6221__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_7111_)
);

FILL FILL_0__16802_ (
);

FILL FILL_0__19274_ (
);

FILL FILL252320x34580 (
);

FILL FILL_0__9375_ (
);

OR2X2 _11646_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_1649_)
);

OR2X2 _11226_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_1429_)
);

FILL FILL427120x44460 (
);

FILL FILL_0__12722_ (
);

FILL FILL162640x69160 (
);

FILL FILL317680x64220 (
);

FILL FILL341240x281580 (
);

FILL FILL_0__15194_ (
);

FILL FILL47880x93860 (
);

FILL FILL433200x237120 (
);

FILL FILL258400x291460 (
);

FILL FILL_0__13507_ (
);

FILL FILL463600x34580 (
);

AND2X2 _16684_ (
    .A(_4214__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_5620_)
);

OR2X2 _16264_ (
    .A(_5202_),
    .B(_5205_),
    .Y(_5206_)
);

FILL FILL_1__9536_ (
);

FILL FILL38760x202540 (
);

FILL FILL256120x34580 (
);

FILL FILL_0__17760_ (
);

FILL FILL_1__10854_ (
);

FILL FILL395200x217360 (
);

FILL FILL166440x69160 (
);

OR2X2 _17889_ (
    .A(_6806_),
    .B(_6805_),
    .Y(_6807_)
);

OR2X2 _17469_ (
    .A(_6393_),
    .B(_6392_),
    .Y(_6394_)
);

OR2X2 _17049_ (
    .A(_5963_),
    .B(_5978_),
    .Y(_5979_)
);

DFFSR _12184_ (
    .CLK(clk_bF$buf80),
    .D(_1851_[19]),
    .Q(\datapath_1.regfile_1.regOut[29] [19]),
    .R(rst_bF$buf76),
    .S(vdd)
);

FILL FILL_0__18965_ (
);

FILL FILL55480x118560 (
);

AND2X2 _18830_ (
    .A(_6297__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_7734_)
);

FILL FILL_0__18125_ (
);

AND2X2 _18410_ (
    .A(_6232__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_7320_)
);

FILL FILL95000x227240 (
);

FILL FILL_0__13680_ (
);

FILL FILL_0__13260_ (
);

FILL FILL_1__11219_ (
);

FILL FILL_0__8646_ (
);

OR2X2 _10917_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_1263_)
);

FILL FILL72960x128440 (
);

NAND3X1 _13389_ (
    .A(ALUControl[1]),
    .B(\datapath_1.alu_1.ALUInB [3]),
    .C(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2926_)
);

FILL FILL129960x133380 (
);

FILL FILL59280x360620 (
);

DFFSR _14750_ (
    .CLK(clk_bF$buf15),
    .D(_3804_[27]),
    .Q(\datapath_1.a [27]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL_0__14045_ (
);

OR2X2 _14330_ (
    .A(vdd),
    .B(ALUOut[30]),
    .Y(_3666_)
);

FILL FILL152000x326040 (
);

FILL FILL477280x247000 (
);

FILL FILL311600x370500 (
);

OR2X2 _15955_ (
    .A(_4900_),
    .B(_4901_),
    .Y(_4902_)
);

OR2X2 _15535_ (
    .A(_4485_),
    .B(_4488_),
    .Y(_4489_)
);

AND2X2 _15115_ (
    .A(_4059_),
    .B(_4013_),
    .Y(_4094_)
);

AND2X2 _10670_ (
    .A(_1138_),
    .B(_1137_),
    .Y(_1125_[6])
);

DFFSR _10250_ (
    .CLK(clk_bF$buf71),
    .D(_861_[20]),
    .Q(\datapath_1.regfile_1.regOut[14] [20]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL_1__8807_ (
);

FILL FILL_1__12597_ (
);

FILL FILL442320x355680 (
);

FILL FILL_1__18823_ (
);

OR2X2 _11875_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_1784__bF$buf3),
    .Y(_1762_)
);

FILL FILL_0__9184_ (
);

OR2X2 _11455_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .B(_1586__bF$buf4),
    .Y(_1542_)
);

DFFSR _11035_ (
    .CLK(clk_bF$buf57),
    .D(_1257_[31]),
    .Q(\datapath_1.regfile_1.regOut[20] [31]),
    .R(rst_bF$buf81),
    .S(vdd)
);

FILL FILL28880x291460 (
);

FILL FILL_0__17816_ (
);

FILL FILL_0__12531_ (
);

FILL FILL491720x153140 (
);

FILL FILL_0__12111_ (
);

FILL FILL254600x187720 (
);

DFFSR _9603_ (
    .CLK(clk_bF$buf22),
    .D(_531_[18]),
    .Q(\datapath_1.regfile_1.regOut[9] [18]),
    .R(rst_bF$buf74),
    .S(vdd)
);

FILL FILL_0__13736_ (
);

AND2X2 _13601_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [1]),
    .Y(_3095_)
);

AND2X2 _16493_ (
    .A(_4208__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_5432_)
);

OR2X2 _16073_ (
    .A(_5017_),
    .B(_5010_),
    .Y(_5018_)
);

FILL FILL_1__15528_ (
);

FILL FILL_1__10663_ (
);

AND2X2 _14806_ (
    .A(_3903_),
    .B(_3902_),
    .Y(_3870_[16])
);

FILL FILL356440x49400 (
);

OR2X2 _17698_ (
    .A(_6615_),
    .B(_6618_),
    .Y(_6619_)
);

AND2X2 _17278_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_6204_)
);

FILL FILL_0__18774_ (
);

FILL FILL_0__18354_ (
);

FILL FILL353400x306280 (
);

FILL FILL239400x330980 (
);

FILL FILL22800x98800 (
);

FILL FILL_0__8875_ (
);

FILL FILL_0__8455_ (
);

OR2X2 _10726_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .B(_1190__bF$buf3),
    .Y(_1176_)
);

OR2X2 _10306_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .B(_992__bF$buf2),
    .Y(_956_)
);

FILL FILL405840x59280 (
);

OR2X2 _13198_ (
    .A(_2212_),
    .B(_2746_),
    .Y(_2747_)
);

FILL FILL_0__19559_ (
);

OR2X2 _19424_ (
    .A(_8285_),
    .B(_8318_),
    .Y(_8319_)
);

FILL FILL_0__19139_ (
);

AND2X2 _19004_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_7905_)
);

FILL FILL_0__14694_ (
);

FILL FILL243960x247000 (
);

FILL FILL179360x326040 (
);

FILL FILL_1__16486_ (
);

AND2X2 _15764_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_4714_)
);

FILL FILL_0__15479_ (
);

FILL FILL_0__15059_ (
);

AND2X2 _15344_ (
    .A(_4167__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_4301_)
);

FILL FILL5320x138320 (
);

FILL FILL165680x350740 (
);

FILL FILL_0__10194_ (
);

FILL FILL_0__16420_ (
);

FILL FILL_0__16000_ (
);

FILL FILL223440x133380 (
);

FILL FILL409640x59280 (
);

OR2X2 _16969_ (
    .A(_5899_),
    .B(_5892_),
    .Y(_5900_)
);

FILL FILL484120x79040 (
);

AND2X2 _16549_ (
    .A(_4197__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_5487_)
);

OR2X2 _16129_ (
    .A(_5069_),
    .B(_5072_),
    .Y(_5073_)
);

AND2X2 _11684_ (
    .A(_1654_),
    .B(_1717_),
    .Y(_1653_[0])
);

FILL FILL461320x335920 (
);

DFFSR _11264_ (
    .CLK(clk_bF$buf56),
    .D(_1389_[2]),
    .Q(\datapath_1.regfile_1.regOut[22] [2]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL_0__17625_ (
);

OR2X2 _17910_ (
    .A(_6827_),
    .B(_6824_),
    .Y(_6828_)
);

FILL FILL_0__12760_ (
);

FILL FILL_0__12340_ (
);

FILL FILL402040x321100 (
);

OR2X2 _9832_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .B(_728__bF$buf4),
    .Y(_720_)
);

OR2X2 _9412_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .B(_530__bF$buf1),
    .Y(_500_)
);

NAND3X1 _12889_ (
    .A(_2453_),
    .B(_2288_),
    .C(_2280_),
    .Y(_2454_)
);

AND2X2 _12469_ (
    .A(_2059_),
    .B(_2061_),
    .Y(_2062_)
);

DFFSR _12049_ (
    .CLK(clk_bF$buf85),
    .D(_1785_[13]),
    .Q(\datapath_1.regfile_1.regOut[28] [13]),
    .R(rst_bF$buf109),
    .S(vdd)
);

FILL FILL_1__14972_ (
);

FILL FILL_0__13965_ (
);

AND2X2 _13830_ (
    .A(_3286_),
    .B(_3285_),
    .Y(\datapath_1.alu_1.ALUInA [4])
);

FILL FILL_0__13545_ (
);

FILL FILL_0__13125_ (
);

XOR2X1 _13410_ (
    .A(_2182_),
    .B(_2391_),
    .Y(_2946_)
);

FILL FILL_1__9574_ (
);

FILL FILL_1__10472_ (
);

DFFSR _14615_ (
    .CLK(clk_bF$buf40),
    .D(_3738_[21]),
    .Q(\datapath_1.PCJump [23]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL500080x167960 (
);

AND2X2 _17087_ (
    .A(_4151__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_6016_)
);

FILL FILL_1__19170_ (
);

AND2X2 _10955_ (
    .A(_1288_),
    .B(_1287_),
    .Y(_1257_[15])
);

AND2X2 _10535_ (
    .A(_1068_),
    .B(_1067_),
    .Y(_1059_[4])
);

DFFSR _10115_ (
    .CLK(clk_bF$buf3),
    .D(_795_[14]),
    .Q(\datapath_1.regfile_1.regOut[13] [14]),
    .R(rst_bF$buf4),
    .S(vdd)
);

FILL FILL91200x93860 (
);

FILL FILL9880x9880 (
);

FILL FILL_0__11611_ (
);

FILL FILL_0__19368_ (
);

OR2X2 _19233_ (
    .A(_8129_),
    .B(_8128_),
    .Y(_8130_)
);

FILL FILL_0__14083_ (
);

FILL FILL_0__9889_ (
);

FILL FILL_1__13403_ (
);

OR2X2 _15993_ (
    .A(_4908_),
    .B(_4939_),
    .Y(_4940_)
);

AND2X2 _15573_ (
    .A(_4241__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_4526_)
);

AND2X2 _15153_ (
    .A(_4112_),
    .B(_4011_),
    .Y(_4118_)
);

FILL FILL24320x217360 (
);

FILL FILL328320x128440 (
);

FILL FILL373160x232180 (
);

FILL FILL301720x9880 (
);

AND2X2 _16778_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_5712_)
);

OR2X2 _16358_ (
    .A(_5297_),
    .B(_5298_),
    .Y(_5299_)
);

OR2X2 _11493_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_1567_)
);

OR2X2 _11073_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_1347_)
);

FILL FILL_0__17854_ (
);

FILL FILL_0__17434_ (
);

FILL FILL_0__17014_ (
);

AND2X2 _9641_ (
    .A(_612_),
    .B(_611_),
    .Y(_597_[7])
);

DFFSR _9221_ (
    .CLK(clk_bF$buf87),
    .D(_333_[23]),
    .Q(\datapath_1.regfile_1.regOut[6] [23]),
    .R(rst_bF$buf54),
    .S(vdd)
);

FILL FILL345040x365560 (
);

NAND2X1 _12698_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2263_)
);

AND2X2 _12278_ (
    .A(_1970_),
    .B(_1969_),
    .Y(_1917_[26])
);

OR2X2 _18924_ (
    .A(_7824_),
    .B(_7825_),
    .Y(_7826_)
);

FILL FILL377720x113620 (
);

FILL FILL_0__18219_ (
);

AND2X2 _18504_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_7413_)
);

FILL FILL_0__13354_ (
);

FILL FILL_1__9383_ (
);

FILL FILL102600x247000 (
);

FILL FILL193040x276640 (
);

FILL FILL_1__15986_ (
);

FILL FILL_1__10281_ (
);

FILL FILL16720x232180 (
);

FILL FILL_0__14979_ (
);

OR2X2 _14844_ (
    .A(\datapath_1.rd2 [29]),
    .B(_3935__bF$buf0),
    .Y(_3929_)
);

FILL FILL_0__14559_ (
);

OR2X2 _14424_ (
    .A(memoryOutData[18]),
    .B(_3737__bF$buf2),
    .Y(_3709_)
);

OR2X2 _14004_ (
    .A(_3421_),
    .B(_3422_),
    .Y(_3423_)
);

FILL FILL117800x14820 (
);

FILL FILL202920x340860 (
);

FILL FILL275880x29640 (
);

FILL FILL_0__15920_ (
);

FILL FILL_0__15500_ (
);

FILL FILL_0__18392_ (
);

FILL FILL345040x59280 (
);

FILL FILL392920x197600 (
);

AND2X2 _15629_ (
    .A(_4230__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_4581_)
);

AND2X2 _15209_ (
    .A(_4166_),
    .B(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_4167_)
);

DFFSR _10764_ (
    .CLK(clk_bF$buf110),
    .D(_1125_[18]),
    .Q(\datapath_1.regfile_1.regOut[18] [18]),
    .R(rst_bF$buf74),
    .S(vdd)
);

FILL FILL_0__10479_ (
);

OR2X2 _10344_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_981_)
);

FILL FILL_0__11000_ (
);

AND2X2 _19462_ (
    .A(_8343_),
    .B(_8342_),
    .Y(_8320_[11])
);

OR2X2 _19042_ (
    .A(_7941_),
    .B(_7938_),
    .Y(_7942_)
);

AND2X2 _8912_ (
    .A(_246_),
    .B(_245_),
    .Y(_201_[22])
);

FILL FILL_0__9698_ (
);

AND2X2 _11969_ (
    .A(_1804_),
    .B(_1803_),
    .Y(_1785_[9])
);

FILL FILL_0__9278_ (
);

DFFSR _11549_ (
    .CLK(clk_bF$buf88),
    .D(_1521_[29]),
    .Q(\datapath_1.regfile_1.regOut[24] [29]),
    .R(rst_bF$buf95),
    .S(vdd)
);

AND2X2 _11129_ (
    .A(_1384_),
    .B(_1383_),
    .Y(_1323_[30])
);

FILL FILL279680x29640 (
);

AND2X2 _12910_ (
    .A(_2456_),
    .B(_2474_),
    .Y(_2475_)
);

FILL FILL_0__12625_ (
);

FILL FILL424840x251940 (
);

FILL FILL_1_BUFX2_insert407 (
);

FILL FILL_1_BUFX2_insert409 (
);

FILL FILL_0__15097_ (
);

OR2X2 _15382_ (
    .A(_4337_),
    .B(_4336_),
    .Y(_4338_)
);

FILL FILL37240x256880 (
);

FILL FILL199880x44460 (
);

FILL FILL_1__14417_ (
);

AND2X2 _16587_ (
    .A(_4223__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_5524_)
);

OR2X2 _16167_ (
    .A(_5107_),
    .B(_5110_),
    .Y(_5111_)
);

FILL FILL_1__18250_ (
);

FILL FILL478040x227240 (
);

FILL FILL_0__17243_ (
);

DFFSR _9870_ (
    .CLK(clk_bF$buf36),
    .D(_663_[27]),
    .Q(\datapath_1.regfile_1.regOut[11] [27]),
    .R(rst_bF$buf78),
    .S(vdd)
);

OR2X2 _9450_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_525_)
);

OR2X2 _9030_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_305_)
);

FILL FILL_1__19035_ (
);

OR2X2 _12087_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_1863_)
);

FILL FILL_0__18868_ (
);

AND2X2 _18733_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_7638_)
);

FILL FILL_0__18448_ (
);

AND2X2 _18313_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_7225_)
);

FILL FILL_0__13583_ (
);

FILL FILL_0__13163_ (
);

FILL FILL504640x207480 (
);

FILL FILL_0__8549_ (
);

FILL FILL_1__12903_ (
);

FILL FILL304760x98800 (
);

OR2X2 _19518_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8381_)
);

FILL FILL_0__14788_ (
);

AND2X2 _14653_ (
    .A(_3821_),
    .B(_3820_),
    .Y(_3804_[8])
);

FILL FILL_0__14368_ (
);

OR2X2 _14233_ (
    .A(MemToReg_bF$buf0),
    .B(ALUOut[30]),
    .Y(_3600_)
);

FILL FILL275120x0 (
);

FILL FILL147440x261820 (
);

OR2X2 _15858_ (
    .A(_4805_),
    .B(_4806_),
    .Y(_4807_)
);

FILL FILL284240x321100 (
);

AND2X2 _15438_ (
    .A(_4154__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_4393_)
);

NOR3X1 _15018_ (
    .A(_4006_),
    .B(_4005_),
    .C(\datapath_1.a3 [2]),
    .Y(_4007_)
);

OR2X2 _10993_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .B(_1322__bF$buf0),
    .Y(_1314_)
);

FILL FILL_1__17941_ (
);

FILL FILL234080x172900 (
);

FILL FILL_0__10288_ (
);

OR2X2 _10573_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .B(_1124__bF$buf1),
    .Y(_1094_)
);

OR2X2 _10153_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .B(_926__bF$buf3),
    .Y(_874_)
);

FILL FILL_0__16934_ (
);

FILL FILL_0__16514_ (
);

FILL FILL33440x286520 (
);

OR2X2 _19271_ (
    .A(_8167_),
    .B(_8166_),
    .Y(_8168_)
);

FILL FILL447640x0 (
);

OR2X2 _8721_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_139_)
);

DFFSR _11778_ (
    .CLK(clk_bF$buf105),
    .D(_1653_[0]),
    .Q(\datapath_1.regfile_1.regOut[26] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

OR2X2 _11358_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_1497_)
);

FILL FILL181640x187720 (
);

FILL FILL_1__13021_ (
);

FILL FILL_0__17719_ (
);

FILL FILL_0__12854_ (
);

FILL FILL_0__12014_ (
);

OR2X2 _15191_ (
    .A(_4137_),
    .B(_4148_),
    .Y(_4149_)
);

AND2X2 _9926_ (
    .A(_762_),
    .B(_761_),
    .Y(_729_[16])
);

AND2X2 _9506_ (
    .A(_542_),
    .B(_541_),
    .Y(_531_[5])
);

FILL FILL369360x172900 (
);

FILL FILL_1__14226_ (
);

FILL FILL308560x281580 (
);

FILL FILL299440x177840 (
);

OR2X2 _13924_ (
    .A(_3354_),
    .B(_3349_),
    .Y(\datapath_1.alu_1.ALUInB [0])
);

FILL FILL_0__13219_ (
);

OR2X2 _13504_ (
    .A(IorD_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [5]),
    .Y(_3024_)
);

OR2X2 _16396_ (
    .A(_5334_),
    .B(_5335_),
    .Y(_5336_)
);

FILL FILL253080x158080 (
);

FILL FILL_1__9668_ (
);

FILL FILL167200x83980 (
);

FILL FILL_0__17892_ (
);

FILL FILL_0__17472_ (
);

FILL FILL228000x24700 (
);

OR2X2 _14709_ (
    .A(\datapath_1.rd1 [27]),
    .B(_3869__bF$buf3),
    .Y(_3859_)
);

FILL FILL_1_CLKBUF1_insert113 (
);

FILL FILL_1_CLKBUF1_insert115 (
);

FILL FILL_1_CLKBUF1_insert117 (
);

FILL FILL_1__19264_ (
);

AND2X2 _18962_ (
    .A(_6323__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_7864_)
);

OR2X2 _18542_ (
    .A(_7449_),
    .B(_7448_),
    .Y(_7450_)
);

FILL FILL_0__18257_ (
);

OR2X2 _18122_ (
    .A(_7021_),
    .B(_7036_),
    .Y(_7037_)
);

FILL FILL268280x4940 (
);

FILL FILL449920x222300 (
);

FILL FILL_0__8778_ (
);

FILL FILL25840x167960 (
);

DFFSR _10629_ (
    .CLK(clk_bF$buf75),
    .D(_1059_[12]),
    .Q(\datapath_1.regfile_1.regOut[17] [12]),
    .R(rst_bF$buf27),
    .S(vdd)
);

OR2X2 _10209_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_911_)
);

FILL FILL388360x158080 (
);

FILL FILL242440x74100 (
);

FILL FILL_0__11705_ (
);

FILL FILL504640x345800 (
);

AND2X2 _19327_ (
    .A(_6271__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_8223_)
);

DFFSR _14882_ (
    .CLK(clk_bF$buf98),
    .D(_3870_[30]),
    .Q(_2_[30]),
    .R(rst_bF$buf61),
    .S(vdd)
);

FILL FILL_0__14177_ (
);

OR2X2 _14462_ (
    .A(vdd),
    .B(\datapath_1.Data [31]),
    .Y(_3734_)
);

OR2X2 _14042_ (
    .A(_3455_),
    .B(_3454_),
    .Y(_3456_)
);

FILL FILL119320x326040 (
);

AND2X2 _15667_ (
    .A(_4142__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_4619_)
);

OR2X2 _15247_ (
    .A(_4201_),
    .B(_4204_),
    .Y(_4205_)
);

FILL FILL269800x74100 (
);

FILL FILL105640x350740 (
);

DFFSR _10382_ (
    .CLK(clk_bF$buf45),
    .D(_927_[23]),
    .Q(\datapath_1.regfile_1.regOut[15] [23]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL470440x24700 (
);

FILL FILL200640x59280 (
);

FILL FILL_0__16743_ (
);

FILL FILL_0__16323_ (
);

OR2X2 _19080_ (
    .A(_7979_),
    .B(_7976_),
    .Y(_7980_)
);

DFFSR _8950_ (
    .CLK(clk_bF$buf33),
    .D(_201_[10]),
    .Q(\datapath_1.regfile_1.regOut[4] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

OR2X2 _8530_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_68__bF$buf4),
    .Y(_52_)
);

FILL FILL427120x182780 (
);

FILL FILL109440x271700 (
);

OR2X2 _11587_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .B(_1652__bF$buf3),
    .Y(_1610_)
);

FILL FILL_1__18115_ (
);

OR2X2 _11167_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(_1454__bF$buf4),
    .Y(_1390_)
);

FILL FILL_0__17948_ (
);

AND2X2 _17813_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_6732_)
);

FILL FILL_0__17108_ (
);

FILL FILL444600x192660 (
);

FILL FILL_0__12663_ (
);

FILL FILL_0__12243_ (
);

FILL FILL409640x355680 (
);

DFFSR _9735_ (
    .CLK(clk_bF$buf1),
    .D(_597_[21]),
    .Q(\datapath_1.regfile_1.regOut[10] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

OR2X2 _9315_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_455_)
);

FILL FILL419520x19760 (
);

FILL FILL_0__13448_ (
);

OR2X2 _13733_ (
    .A(_3206_),
    .B(_3207_),
    .Y(_3208_)
);

FILL FILL_0__13028_ (
);

OR2X2 _13313_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .B(_2853_),
    .Y(_2854_)
);

FILL FILL494000x39520 (
);

AND2X2 _14938_ (
    .A(_3971_),
    .B(_3970_),
    .Y(_3936_[17])
);

AND2X2 _14518_ (
    .A(_3751_),
    .B(_3750_),
    .Y(_3738_[6])
);

FILL FILL316160x34580 (
);

OR2X2 _18771_ (
    .A(_7675_),
    .B(_7668_),
    .Y(_7676_)
);

FILL FILL_0__18486_ (
);

FILL FILL_0__18066_ (
);

AND2X2 _18351_ (
    .A(_6282__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_7262_)
);

FILL FILL_0__8587_ (
);

OR2X2 _10858_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .B(_1256__bF$buf0),
    .Y(_1244_)
);

OR2X2 _10438_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .B(_1058__bF$buf0),
    .Y(_1024_)
);

OR2X2 _10018_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .B(_860__bF$buf1),
    .Y(_804_)
);

FILL FILL_1__12101_ (
);

FILL FILL215840x128440 (
);

FILL FILL_0__11514_ (
);

AND2X2 _19556_ (
    .A(_8386_),
    .B(BranchNe),
    .Y(_8387_)
);

OR2X2 _19136_ (
    .A(_8034_),
    .B(_8033_),
    .Y(_8035_)
);

OR2X2 _14691_ (
    .A(\datapath_1.rd1 [21]),
    .B(_3869__bF$buf1),
    .Y(_3847_)
);

OR2X2 _14271_ (
    .A(\datapath_1.ALUResult [10]),
    .B(_3671__bF$buf2),
    .Y(_3627_)
);

FILL FILL479560x177840 (
);

FILL FILL93480x172900 (
);

FILL FILL_0__12719_ (
);

OR2X2 _15896_ (
    .A(_4843_),
    .B(_4836_),
    .Y(_4844_)
);

AND2X2 _15476_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_4431_)
);

AND2X2 _15056_ (
    .A(_4022_),
    .B(RegWrite),
    .Y(_4045_)
);

OR2X2 _10191_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_899_)
);

FILL FILL_0__16972_ (
);

FILL FILL_0__16552_ (
);

FILL FILL310840x345800 (
);

FILL FILL150480x271700 (
);

FILL FILL374680x34580 (
);

FILL FILL456760x202540 (
);

FILL FILL236360x286520 (
);

FILL FILL_1__18764_ (
);

FILL FILL72200x256880 (
);

DFFSR _11396_ (
    .CLK(clk_bF$buf68),
    .D(_1455_[5]),
    .Q(\datapath_1.regfile_1.regOut[23] [5]),
    .R(rst_bF$buf21),
    .S(vdd)
);

FILL FILL69160x207480 (
);

AND2X2 _17622_ (
    .A(_6262__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_6544_)
);

FILL FILL_0__17337_ (
);

OR2X2 _17202_ (
    .A(_6128_),
    .B(_6129_),
    .Y(_6130_)
);

FILL FILL376200x167960 (
);

FILL FILL_0__12472_ (
);

FILL FILL463600x172900 (
);

FILL FILL428640x335920 (
);

OR2X2 _9964_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .B(_794__bF$buf3),
    .Y(_788_)
);

OR2X2 _9544_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .B(_596__bF$buf2),
    .Y(_568_)
);

OR2X2 _9124_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .B(_398__bF$buf1),
    .Y(_348_)
);

FILL FILL_1__19129_ (
);

FILL FILL107920x237120 (
);

FILL FILL505400x79040 (
);

OR2X2 _18827_ (
    .A(_7730_),
    .B(_7729_),
    .Y(_7731_)
);

FILL FILL_0_BUFX2_insert440 (
);

FILL FILL198360x266760 (
);

FILL FILL412680x49400 (
);

FILL FILL_0_BUFX2_insert441 (
);

AND2X2 _18407_ (
    .A(_6247__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_7317_)
);

FILL FILL126160x306280 (
);

FILL FILL_0_BUFX2_insert443 (
);

OR2X2 _13962_ (
    .A(_3385_),
    .B(_3386_),
    .Y(_3387_)
);

FILL FILL_0__13677_ (
);

FILL FILL213560x311220 (
);

FILL FILL_0_BUFX2_insert445 (
);

AND2X2 _13542_ (
    .A(_3049_),
    .B(_3048_),
    .Y(_1_[17])
);

NAND2X1 _13122_ (
    .A(_2674_),
    .B(_2672_),
    .Y(_2675_)
);

FILL FILL_0_BUFX2_insert447 (
);

FILL FILL_0_BUFX2_insert449 (
);

FILL FILL_1__9286_ (
);

FILL FILL143640x316160 (
);

FILL FILL_0__17090_ (
);

FILL FILL133000x276640 (
);

FILL FILL_1__15469_ (
);

DFFSR _14747_ (
    .CLK(clk_bF$buf41),
    .D(_3804_[24]),
    .Q(\datapath_1.a [24]),
    .R(rst_bF$buf63),
    .S(vdd)
);

OR2X2 _14327_ (
    .A(vdd),
    .B(ALUOut[29]),
    .Y(_3664_)
);

FILL FILL_1__16410_ (
);

FILL FILL110960x177840 (
);

FILL FILL_0__15403_ (
);

FILL FILL357200x113620 (
);

FILL FILL_0__18295_ (
);

AND2X2 _18580_ (
    .A(_7487_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.rd1 [18])
);

AND2X2 _18160_ (
    .A(_6297__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_7074_)
);

FILL FILL416480x49400 (
);

FILL FILL503880x340860 (
);

FILL FILL368600x182780 (
);

FILL FILL_0__8396_ (
);

FILL FILL_1__17615_ (
);

AND2X2 _10667_ (
    .A(_1136_),
    .B(_1135_),
    .Y(_1125_[5])
);

DFFSR _10247_ (
    .CLK(clk_bF$buf8),
    .D(_861_[17]),
    .Q(\datapath_1.regfile_1.regOut[14] [17]),
    .R(rst_bF$buf10),
    .S(vdd)
);

FILL FILL_0__16608_ (
);

FILL FILL_0__11743_ (
);

FILL FILL_0__11323_ (
);

AND2X2 _19365_ (
    .A(_6289__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_8260_)
);

AND2X2 _14080_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3488_)
);

DFFSR _8815_ (
    .CLK(clk_bF$buf45),
    .D(_135_[4]),
    .Q(\datapath_1.regfile_1.regOut[3] [4]),
    .R(rst_bF$buf54),
    .S(vdd)
);

FILL FILL351880x251940 (
);

FILL FILL65360x237120 (
);

FILL FILL_0__12948_ (
);

FILL FILL388360x311220 (
);

OR2X2 _12813_ (
    .A(gnd),
    .B(ALUControl[2]),
    .Y(_2378_)
);

FILL FILL_0__12108_ (
);

FILL FILL125400x291460 (
);

OR2X2 _15285_ (
    .A(_4240_),
    .B(_4242_),
    .Y(_4243_)
);

FILL FILL482600x34580 (
);

FILL FILL_1__8977_ (
);

FILL FILL_0__16361_ (
);

FILL FILL185440x69160 (
);

FILL FILL209760x113620 (
);

FILL FILL_0__17986_ (
);

FILL FILL_0__17566_ (
);

AND2X2 _17851_ (
    .A(_6289__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_6770_)
);

OR2X2 _17431_ (
    .A(_6351_),
    .B(_6355_),
    .Y(_6356_)
);

AND2X2 _17011_ (
    .A(_4228__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_5942_)
);

FILL FILL343520x281580 (
);

FILL FILL262200x217360 (
);

FILL FILL386840x345800 (
);

AND2X2 _9773_ (
    .A(_680_),
    .B(_679_),
    .Y(_663_[8])
);

DFFSR _9353_ (
    .CLK(clk_bF$buf55),
    .D(_399_[26]),
    .Q(\datapath_1.regfile_1.regOut[7] [26]),
    .R(rst_bF$buf14),
    .S(vdd)
);

OR2X2 _18636_ (
    .A(_7542_),
    .B(_7541_),
    .Y(_7543_)
);

OR2X2 _18216_ (
    .A(_7128_),
    .B(_7127_),
    .Y(_7129_)
);

FILL FILL226480x350740 (
);

OR2X2 _13771_ (
    .A(_3240_),
    .B(_3239_),
    .Y(_3241_)
);

FILL FILL_0__13066_ (
);

OAI21X1 _13351_ (
    .A(_2402_),
    .B(_2185_),
    .C(_2198_),
    .Y(_2890_)
);

FILL FILL_0__9813_ (
);

FILL FILL189240x69160 (
);

OR2X2 _14976_ (
    .A(\datapath_1.mux_pcsrc.dout [30]),
    .B(_4001__bF$buf4),
    .Y(_3997_)
);

OR2X2 _14556_ (
    .A(memoryOutData[19]),
    .B(_3803__bF$buf2),
    .Y(_3777_)
);

AND2X2 _14136_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3536_)
);

FILL FILL_0__15632_ (
);

FILL FILL_0__15212_ (
);

FILL FILL254600x232180 (
);

DFFSR _10896_ (
    .CLK(clk_bF$buf98),
    .D(_1191_[21]),
    .Q(\datapath_1.regfile_1.regOut[19] [21]),
    .R(rst_bF$buf87),
    .S(vdd)
);

OR2X2 _10476_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_1049_)
);

OR2X2 _10056_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_829_)
);

FILL FILL_0__16837_ (
);

AND2X2 _16702_ (
    .A(_4214__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_5637_)
);

FILL FILL_0__16417_ (
);

FILL FILL_0__11552_ (
);

FILL FILL_0__11132_ (
);

AND2X2 _19174_ (
    .A(_6328__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_8072_)
);

AND2X2 _8624_ (
    .A(_94_),
    .B(_93_),
    .Y(_69_[12])
);

FILL FILL_1__18629_ (
);

FILL FILL_1__13344_ (
);

AND2X2 _17907_ (
    .A(_6255__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_6825_)
);

XNOR2X1 _12622_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2187_)
);

OR2X2 _12202_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .B(_1982__bF$buf2),
    .Y(_1920_)
);

AND2X2 _15094_ (
    .A(_4041_),
    .B(_4077_),
    .Y(_4078_)
);

FILL FILL273600x54340 (
);

OR2X2 _9829_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .B(_728__bF$buf2),
    .Y(_718_)
);

OR2X2 _9409_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .B(_530__bF$buf1),
    .Y(_498_)
);

FILL FILL_0__16590_ (
);

FILL FILL41040x340860 (
);

AND2X2 _13827_ (
    .A(_3284_),
    .B(_3283_),
    .Y(\datapath_1.alu_1.ALUInA [3])
);

OR2X2 _13407_ (
    .A(_2498_),
    .B(_2929_),
    .Y(_2943_)
);

FILL FILL_1__15910_ (
);

OR2X2 _16299_ (
    .A(_5240_),
    .B(_5239_),
    .Y(_5241_)
);

FILL FILL_0__14903_ (
);

FILL FILL_1__18382_ (
);

FILL FILL55480x301340 (
);

FILL FILL180880x118560 (
);

AND2X2 _17660_ (
    .A(_6328__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_6582_)
);

FILL FILL_0__17375_ (
);

OR2X2 _17240_ (
    .A(_6166_),
    .B(_6159_),
    .Y(_6167_)
);

FILL FILL448400x276640 (
);

FILL FILL_1__10049_ (
);

FILL FILL76000x247000 (
);

FILL FILL399000x321100 (
);

OR2X2 _9582_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_593_)
);

OR2X2 _9162_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_373_)
);

FILL FILL62320x271700 (
);

FILL FILL289560x217360 (
);

FILL FILL442320x88920 (
);

FILL FILL_0__10823_ (
);

FILL FILL_0__10403_ (
);

AND2X2 _18865_ (
    .A(_6264__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_7768_)
);

FILL FILL_0_BUFX2_insert820 (
);

FILL FILL_0_BUFX2_insert821 (
);

OR2X2 _18445_ (
    .A(_7354_),
    .B(_7351_),
    .Y(_7355_)
);

AND2X2 _18025_ (
    .A(_6282__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_6941_)
);

FILL FILL_0_BUFX2_insert823 (
);

FILL FILL_0__13295_ (
);

OR2X2 _13580_ (
    .A(ALUOut[30]),
    .B(_3079__bF$buf3),
    .Y(_3075_)
);

FILL FILL_0_BUFX2_insert825 (
);

NAND3X1 _13160_ (
    .A(_2666_),
    .B(_2293_),
    .C(_2524_),
    .Y(_2711_)
);

FILL FILL_0_BUFX2_insert827 (
);

FILL FILL_0_BUFX2_insert829 (
);

FILL FILL_0__19521_ (
);

FILL FILL_0__19101_ (
);

FILL FILL_0__9622_ (
);

FILL FILL_1__15087_ (
);

AND2X2 _14785_ (
    .A(_3889_),
    .B(_3888_),
    .Y(_3870_[9])
);

DFFSR _14365_ (
    .CLK(clk_bF$buf20),
    .D(_3606_[29]),
    .Q(ALUOut[29]),
    .R(rst_bF$buf91),
    .S(vdd)
);

FILL FILL497040x167960 (
);

FILL FILL_0__15861_ (
);

FILL FILL_0__15441_ (
);

FILL FILL_0__15021_ (
);

FILL FILL9880x167960 (
);

FILL FILL408880x44460 (
);

FILL FILL82840x74100 (
);

FILL FILL446120x88920 (
);

FILL FILL442320x217360 (
);

FILL FILL_1__17233_ (
);

OR2X2 _10285_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .B(_992__bF$buf4),
    .Y(_942_)
);

OR2X2 _16931_ (
    .A(_5862_),
    .B(_5861_),
    .Y(_5863_)
);

FILL FILL127680x256880 (
);

AND2X2 _16511_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_5449_)
);

FILL FILL254600x370500 (
);

OR2X2 _8853_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_207_)
);

FILL FILL351880x321100 (
);

BUFX2 _8433_ (
    .A(_2_[9]),
    .Y(memoryWriteData[9])
);

FILL FILL_1__13993_ (
);

FILL FILL_1__13573_ (
);

OR2X2 _17716_ (
    .A(_6629_),
    .B(_6636_),
    .Y(_6637_)
);

NAND2X1 _12851_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2416_)
);

FILL FILL_0__12566_ (
);

FILL FILL7600x138320 (
);

DFFSR _12431_ (
    .CLK(clk_bF$buf67),
    .D(_1983_[8]),
    .Q(\datapath_1.regfile_1.regOut[31] [8]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL_0__12146_ (
);

AND2X2 _12011_ (
    .A(_1832_),
    .B(_1831_),
    .Y(_1785_[23])
);

AND2X2 _9638_ (
    .A(_610_),
    .B(_609_),
    .Y(_597_[6])
);

DFFSR _9218_ (
    .CLK(clk_bF$buf56),
    .D(_333_[20]),
    .Q(\datapath_1.regfile_1.regOut[6] [20]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL294120x370500 (
);

FILL FILL_1__14778_ (
);

AND2X2 _13636_ (
    .A(_3087__bF$buf2),
    .B(\datapath_1.ALUResult [6]),
    .Y(_3125_)
);

INVX1 _13216_ (
    .A(_2763_),
    .Y(\datapath_1.ALUResult [14])
);

FILL FILL_0__14712_ (
);

FILL FILL130720x34580 (
);

FILL FILL_0__17184_ (
);

FILL FILL481080x88920 (
);

OR2X2 _9391_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .B(_530__bF$buf1),
    .Y(_486_)
);

FILL FILL_0__15917_ (
);

FILL FILL66880x187720 (
);

FILL FILL161120x9880 (
);

FILL FILL_0__10212_ (
);

FILL FILL215840x79040 (
);

OR2X2 _18674_ (
    .A(_7572_),
    .B(_7579_),
    .Y(_7580_)
);

FILL FILL_0__18389_ (
);

OR2X2 _18254_ (
    .A(_7132_),
    .B(_7166_),
    .Y(_7167_)
);

FILL FILL_1__17709_ (
);

FILL FILL_0__11837_ (
);

FILL FILL_0__9011_ (
);

AND2X2 _11702_ (
    .A(_1666_),
    .B(_1665_),
    .Y(_1653_[6])
);

FILL FILL502360x167960 (
);

AND2X2 _19459_ (
    .A(_8341_),
    .B(_8340_),
    .Y(_8320_[10])
);

AND2X2 _19039_ (
    .A(_6326__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_7939_)
);

DFFSR _14594_ (
    .CLK(clk_bF$buf65),
    .D(_3738_[0]),
    .Q(\aluControl_1.inst [0]),
    .R(rst_bF$buf91),
    .S(vdd)
);

OR2X2 _14174_ (
    .A(\datapath_1.Data [10]),
    .B(_3605__bF$buf0),
    .Y(_3561_)
);

AND2X2 _8909_ (
    .A(_244_),
    .B(_243_),
    .Y(_201_[21])
);

FILL FILL_0__15670_ (
);

FILL FILL146680x370500 (
);

FILL FILL_1__13209_ (
);

FILL FILL_1_BUFX2_insert370 (
);

FILL FILL163400x4940 (
);

AND2X2 _12907_ (
    .A(_2471_),
    .B(_2265_),
    .Y(_2472_)
);

FILL FILL_1_BUFX2_insert372 (
);

FILL FILL_1_BUFX2_insert374 (
);

OR2X2 _15799_ (
    .A(_4748_),
    .B(_4741_),
    .Y(_4749_)
);

OR2X2 _15379_ (
    .A(_4333_),
    .B(_4334_),
    .Y(_4335_)
);

FILL FILL_1__17882_ (
);

AND2X2 _10094_ (
    .A(_854_),
    .B(_853_),
    .Y(_795_[29])
);

AND2X2 _16740_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_5675_)
);

FILL FILL_0__16455_ (
);

FILL FILL_0__16035_ (
);

OR2X2 _16320_ (
    .A(_5260_),
    .B(_5259_),
    .Y(_5261_)
);

FILL FILL_0__11590_ (
);

FILL FILL_0__11170_ (
);

OR2X2 _8662_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .B(_134__bF$buf0),
    .Y(_120_)
);

FILL FILL157320x242060 (
);

FILL FILL340480x44460 (
);

FILL FILL_1__10910_ (
);

OR2X2 _11299_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .B(_1520__bF$buf1),
    .Y(_1458_)
);

OR2X2 _17945_ (
    .A(_6861_),
    .B(_6854_),
    .Y(_6862_)
);

AND2X2 _17525_ (
    .A(_6289__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_6449_)
);

AND2X2 _17105_ (
    .A(_4189__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_6034_)
);

FILL FILL227240x103740 (
);

FILL FILL_0__12795_ (
);

OR2X2 _12660_ (
    .A(_2217_),
    .B(_2224_),
    .Y(_2225_)
);

FILL FILL_0__12375_ (
);

OR2X2 _12240_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_1945_)
);

FILL FILL339720x153140 (
);

FILL FILL_0__18601_ (
);

DFFSR _9867_ (
    .CLK(clk_bF$buf96),
    .D(_663_[24]),
    .Q(\datapath_1.regfile_1.regOut[11] [24]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9447_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_523_)
);

FILL FILL500840x123500 (
);

OR2X2 _9027_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_303_)
);

OR2X2 _13865_ (
    .A(\datapath_1.a [16]),
    .B(_3342__bF$buf2),
    .Y(_3310_)
);

AND2X2 _13445_ (
    .A(_2807_),
    .B(_2778_),
    .Y(_2978_)
);

NAND3X1 _13025_ (
    .A(_2541_),
    .B(_2339_),
    .C(_2524_),
    .Y(_2584_)
);

FILL FILL_0__14941_ (
);

FILL FILL411920x286520 (
);

FILL FILL_0__14521_ (
);

FILL FILL_0__14101_ (
);

FILL FILL75240x242060 (
);

FILL FILL408880x237120 (
);

FILL FILL_0__9907_ (
);

FILL FILL379240x153140 (
);

FILL FILL347320x365560 (
);

FILL FILL_1__16733_ (
);

FILL FILL_0__15726_ (
);

FILL FILL_0__15306_ (
);

FILL FILL364800x375440 (
);

FILL FILL_0__10441_ (
);

FILL FILL196840x34580 (
);

FILL FILL_0__10021_ (
);

AND2X2 _18483_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_7392_)
);

FILL FILL265240x271700 (
);

OR2X2 _18063_ (
    .A(_6976_),
    .B(_6977_),
    .Y(_6978_)
);

FILL FILL195320x276640 (
);

FILL FILL_1__12233_ (
);

FILL FILL_0__9660_ (
);

FILL FILL_0__11646_ (
);

DFFSR _11931_ (
    .CLK(clk_bF$buf6),
    .D(_1719_[24]),
    .Q(\datapath_1.regfile_1.regOut[27] [24]),
    .R(rst_bF$buf31),
    .S(vdd)
);

FILL FILL_0__11226_ (
);

OR2X2 _11511_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_1579_)
);

FILL FILL79040x350740 (
);

OR2X2 _19268_ (
    .A(_8164_),
    .B(_8161_),
    .Y(_8165_)
);

FILL FILL11400x64220 (
);

OR2X2 _8718_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_137_)
);

FILL FILL136800x222300 (
);

FILL FILL483360x261820 (
);

FILL FILL_1__13858_ (
);

FILL FILL_1__13438_ (
);

FILL FILL217360x192660 (
);

INVX1 _12716_ (
    .A(_2280_),
    .Y(_2281_)
);

FILL FILL_1_BUFX2_insert41 (
);

FILL FILL221920x256880 (
);

FILL FILL_1_BUFX2_insert43 (
);

NOR3X1 _15188_ (
    .A(_4145_),
    .B(_4144_),
    .C(_4140_),
    .Y(_4146_)
);

FILL FILL117800x88920 (
);

FILL FILL_0__16684_ (
);

FILL FILL383040x0 (
);

FILL FILL131480x64220 (
);

AND2X2 _8891_ (
    .A(_232_),
    .B(_231_),
    .Y(_201_[15])
);

AND2X2 _8471_ (
    .A(_12_),
    .B(_11_),
    .Y(_3_[4])
);

FILL FILL_1__18056_ (
);

FILL FILL_0__17889_ (
);

AND2X2 _17754_ (
    .A(_6323__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_6674_)
);

FILL FILL_0__17049_ (
);

AND2X2 _17334_ (
    .A(_6259__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_6260_)
);

FILL FILL_0__18830_ (
);

FILL FILL39520x256880 (
);

OR2X2 _9676_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .B(_662__bF$buf3),
    .Y(_636_)
);

OR2X2 _9256_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .B(_464__bF$buf4),
    .Y(_416_)
);

FILL FILL_1__11504_ (
);

FILL FILL_0__8931_ (
);

FILL FILL_0__10917_ (
);

AND2X2 _18959_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_7861_)
);

OR2X2 _18539_ (
    .A(_7446_),
    .B(_7445_),
    .Y(_7447_)
);

OR2X2 _18119_ (
    .A(_7033_),
    .B(_7032_),
    .Y(_7034_)
);

FILL FILL_1_BUFX2_insert1131 (
);

FILL FILL_1_BUFX2_insert1133 (
);

FILL FILL_0__13389_ (
);

OR2X2 _13674_ (
    .A(_3157_),
    .B(_3154_),
    .Y(\datapath_1.mux_pcsrc.dout [11])
);

NAND2X1 _13254_ (
    .A(_2798_),
    .B(_2796_),
    .Y(_2799_)
);

FILL FILL_0__14330_ (
);

FILL FILL289560x83980 (
);

FILL FILL473480x83980 (
);

FILL FILL323000x281580 (
);

DFFSR _14879_ (
    .CLK(clk_bF$buf80),
    .D(_3870_[27]),
    .Q(_2_[27]),
    .R(rst_bF$buf104),
    .S(vdd)
);

OR2X2 _14459_ (
    .A(vdd),
    .B(\datapath_1.Data [30]),
    .Y(_3732_)
);

OR2X2 _14039_ (
    .A(_3451_),
    .B(_3452_),
    .Y(_3453_)
);

FILL FILL505400x192660 (
);

FILL FILL_0__15955_ (
);

FILL FILL_0__15535_ (
);

OR2X2 _15820_ (
    .A(_4768_),
    .B(_4767_),
    .Y(_4769_)
);

OR2X2 _15400_ (
    .A(_4355_),
    .B(_4348_),
    .Y(_4356_)
);

OR2X2 _18292_ (
    .A(_7203_),
    .B(_7202_),
    .Y(_7204_)
);

FILL FILL151240x321100 (
);

FILL FILL346560x133380 (
);

FILL FILL179360x14820 (
);

FILL FILL_1__17747_ (
);

AND2X2 _10799_ (
    .A(_1204_),
    .B(_1203_),
    .Y(_1191_[6])
);

DFFSR _10379_ (
    .CLK(clk_bF$buf100),
    .D(_927_[20]),
    .Q(\datapath_1.regfile_1.regOut[15] [20]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL50160x64220 (
);

FILL FILL46360x143260 (
);

AND2X2 _16605_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_5542_)
);

FILL FILL_0__11875_ (
);

OR2X2 _11740_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .B(_1718__bF$buf2),
    .Y(_1692_)
);

FILL FILL_0__11455_ (
);

FILL FILL449920x158080 (
);

OR2X2 _11320_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .B(_1520__bF$buf1),
    .Y(_1472_)
);

OR2X2 _19497_ (
    .A(gnd),
    .B(_8385__bF$buf2),
    .Y(_8367_)
);

AND2X2 _19077_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_7977_)
);

DFFSR _8947_ (
    .CLK(clk_bF$buf54),
    .D(_201_[7]),
    .Q(\datapath_1.regfile_1.regOut[4] [7]),
    .R(rst_bF$buf48),
    .S(vdd)
);

OR2X2 _8527_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .B(_68__bF$buf0),
    .Y(_50_)
);

FILL FILL149720x261820 (
);

FILL FILL28880x316160 (
);

FILL FILL18240x276640 (
);

FILL FILL_1_BUFX2_insert750 (
);

OR2X2 _12945_ (
    .A(_2387__bF$buf2),
    .B(_2508_),
    .Y(_2509_)
);

FILL FILL_1_BUFX2_insert752 (
);

AND2X2 _12525_ (
    .A(_2112_),
    .B(_2114_),
    .Y(_2115_)
);

OR2X2 _12105_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_1875_)
);

FILL FILL_1_BUFX2_insert754 (
);

FILL FILL236360x172900 (
);

FILL FILL79040x0 (
);

FILL FILL_0__13601_ (
);

FILL FILL358720x360620 (
);

FILL FILL_0__16493_ (
);

FILL FILL_0__16073_ (
);

FILL FILL459040x247000 (
);

FILL FILL186200x83980 (
);

FILL FILL107160x163020 (
);

FILL FILL120080x158080 (
);

FILL FILL86640x103740 (
);

FILL FILL183920x187720 (
);

BUFX2 BUFX2_insert420 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf0 )
);

BUFX2 BUFX2_insert421 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf4)
);

BUFX2 BUFX2_insert422 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf3)
);

BUFX2 BUFX2_insert423 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf2)
);

OR2X2 _17983_ (
    .A(_6899_),
    .B(_6896_),
    .Y(_6900_)
);

BUFX2 BUFX2_insert424 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf1)
);

FILL FILL_0__17698_ (
);

OR2X2 _17563_ (
    .A(_6484_),
    .B(_6485_),
    .Y(_6486_)
);

FILL FILL_0__17278_ (
);

BUFX2 BUFX2_insert425 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf0)
);

BUFX2 BUFX2_insert426 (
    .A(_6221_),
    .Y(_6221__bF$buf4)
);

OR2X2 _17143_ (
    .A(_6064_),
    .B(_6071_),
    .Y(_6072_)
);

BUFX2 BUFX2_insert427 (
    .A(_6221_),
    .Y(_6221__bF$buf3)
);

BUFX2 BUFX2_insert428 (
    .A(_6221_),
    .Y(_6221__bF$buf2)
);

BUFX2 BUFX2_insert429 (
    .A(_6221_),
    .Y(_6221__bF$buf1)
);

FILL FILL12920x311220 (
);

DFFSR _9485_ (
    .CLK(clk_bF$buf0),
    .D(_465_[29]),
    .Q(\datapath_1.regfile_1.regOut[8] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

AND2X2 _9065_ (
    .A(_328_),
    .B(_327_),
    .Y(_267_[30])
);

FILL FILL_1__11313_ (
);

FILL FILL_0__10726_ (
);

AND2X2 _18768_ (
    .A(_6326__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_7673_)
);

OR2X2 _18348_ (
    .A(_7255_),
    .B(_7258_),
    .Y(_7259_)
);

FILL FILL12160x217360 (
);

OR2X2 _13483_ (
    .A(\datapath_1.PCJump [16]),
    .B(_3005_),
    .Y(_3012_)
);

XOR2X1 _13063_ (
    .A(_2267_),
    .B(_2619_),
    .Y(_2620_)
);

FILL FILL_0__19004_ (
);

FILL FILL170240x49400 (
);

FILL FILL_1__12938_ (
);

FILL FILL281200x291460 (
);

FILL FILL_0__9945_ (
);

FILL FILL98800x88920 (
);

FILL FILL_0__9525_ (
);

FILL FILL_0__9105_ (
);

FILL FILL241680x4940 (
);

OR2X2 _14688_ (
    .A(\datapath_1.rd1 [20]),
    .B(_3869__bF$buf1),
    .Y(_3845_)
);

OR2X2 _14268_ (
    .A(\datapath_1.ALUResult [9]),
    .B(_3671__bF$buf4),
    .Y(_3625_)
);

FILL FILL_1__16351_ (
);

OR2X2 _10188_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_897_)
);

FILL FILL_1__12691_ (
);

FILL FILL59280x182780 (
);

FILL FILL_0__16969_ (
);

FILL FILL_0__16549_ (
);

AND2X2 _16834_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_5767_)
);

AND2X2 _16414_ (
    .A(_4241__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_5354_)
);

FILL FILL_0__16129_ (
);

FILL FILL_0__11684_ (
);

AND2X2 _8756_ (
    .A(_162_),
    .B(_161_),
    .Y(_135_[13])
);

OR2X2 _17619_ (
    .A(_6539_),
    .B(_6540_),
    .Y(_6541_)
);

FILL FILL_0__12889_ (
);

NAND2X1 _12754_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2319_)
);

OR2X2 _12334_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .B(_2048__bF$buf1),
    .Y(_1988_)
);

FILL FILL82080x360620 (
);

FILL FILL_0__13830_ (
);

FILL FILL_0__13410_ (
);

FILL FILL63080x197600 (
);

FILL FILL_1__8498_ (
);

OR2X2 _13959_ (
    .A(_3384_),
    .B(_3381_),
    .Y(\datapath_1.alu_1.ALUInB [5])
);

AND2X2 _13539_ (
    .A(_3047_),
    .B(_3046_),
    .Y(_1_[16])
);

MUX2X1 _13119_ (
    .A(_2593_),
    .B(_2548_),
    .S(_2279_),
    .Y(_2672_)
);

FILL FILL_1__15202_ (
);

OR2X2 _14900_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_iord.din0 [5]),
    .Y(_3946_)
);

AND2X2 _17792_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_6712_)
);

AND2X2 _17372_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_6298_)
);

FILL FILL_1__16827_ (
);

OR2X2 _9294_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_441_)
);

FILL FILL_1__11122_ (
);

FILL FILL449160x311220 (
);

FILL FILL_0__10955_ (
);

FILL FILL_0__10535_ (
);

AND2X2 _10820_ (
    .A(_1218_),
    .B(_1217_),
    .Y(_1191_[13])
);

AND2X2 _10400_ (
    .A(_998_),
    .B(_997_),
    .Y(_993_[2])
);

OR2X2 _18997_ (
    .A(_7897_),
    .B(_7894_),
    .Y(_7898_)
);

OR2X2 _18577_ (
    .A(_7469_),
    .B(_7484_),
    .Y(_7485_)
);

AND2X2 _18157_ (
    .A(_6272__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_7071_)
);

AND2X2 _13292_ (
    .A(_2834_),
    .B(_2823_),
    .Y(_2835_)
);

FILL FILL_0__19233_ (
);

FILL FILL497800x98800 (
);

FILL FILL281960x59280 (
);

FILL FILL_0__9754_ (
);

OR2X2 _11605_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_1652__bF$buf4),
    .Y(_1622_)
);

OR2X2 _14497_ (
    .A(\aluControl_1.inst [0]),
    .B(IRWrite_bF$buf0),
    .Y(_3802_)
);

OR2X2 _14077_ (
    .A(_3485_),
    .B(_3484_),
    .Y(_3486_)
);

FILL FILL456760x69160 (
);

FILL FILL_0__15573_ (
);

FILL FILL_0__15153_ (
);

FILL FILL_1__12080_ (
);

FILL FILL_0__16778_ (
);

AND2X2 _16643_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_5579_)
);

FILL FILL_0__16358_ (
);

OR2X2 _16223_ (
    .A(_5165_),
    .B(_5164_),
    .Y(_5166_)
);

FILL FILL_0__11073_ (
);

FILL FILL_1__9915_ (
);

OR2X2 _8985_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_275_)
);

DFFSR _8565_ (
    .CLK(clk_bF$buf28),
    .D(_3_[12]),
    .Q(\datapath_1.regfile_1.regOut[1] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

FILL FILL_1__10813_ (
);

FILL FILL504640x64220 (
);

AND2X2 _17848_ (
    .A(_6271__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [7]),
    .Y(_6767_)
);

INVX1 _17428_ (
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_6353_)
);

AND2X2 _17008_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_5939_)
);

FILL FILL_0__12698_ (
);

AND2X2 _12983_ (
    .A(_2543_),
    .B(_2539_),
    .Y(_2544_)
);

FILL FILL_1__19511_ (
);

FILL FILL_0__12278_ (
);

AND2X2 _12563_ (
    .A(_2083_),
    .B(_2080_),
    .Y(_2084_)
);

AND2X2 _12143_ (
    .A(_1900_),
    .B(_1899_),
    .Y(_1851_[24])
);

FILL FILL261440x9880 (
);

FILL FILL196840x158080 (
);

FILL FILL_0__8605_ (
);

OR2X2 _13768_ (
    .A(_3236_),
    .B(_3237_),
    .Y(_3238_)
);

FILL FILL21280x286520 (
);

AND2X2 _13348_ (
    .A(_2887_),
    .B(_2885_),
    .Y(_2888_)
);

FILL FILL244720x4940 (
);

FILL FILL_1__15851_ (
);

FILL FILL_0__14844_ (
);

BUFX2 BUFX2_insert800 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf2 )
);

BUFX2 BUFX2_insert801 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf1 )
);

BUFX2 BUFX2_insert802 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf0 )
);

BUFX2 BUFX2_insert803 (
    .A(_4177_),
    .Y(_4177__bF$buf4)
);

BUFX2 BUFX2_insert804 (
    .A(_4177_),
    .Y(_4177__bF$buf3)
);

BUFX2 BUFX2_insert805 (
    .A(_4177_),
    .Y(_4177__bF$buf2)
);

BUFX2 BUFX2_insert806 (
    .A(_4177_),
    .Y(_4177__bF$buf1)
);

AND2X2 _17181_ (
    .A(_4217__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_6109_)
);

BUFX2 BUFX2_insert807 (
    .A(_4177_),
    .Y(_4177__bF$buf0)
);

BUFX2 BUFX2_insert808 (
    .A(_6323_),
    .Y(_6323__bF$buf4)
);

BUFX2 BUFX2_insert809 (
    .A(_6323_),
    .Y(_6323__bF$buf3)
);

FILL FILL_1__16216_ (
);

AND2X2 _15914_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_4862_)
);

FILL FILL128440x306280 (
);

FILL FILL_0__10344_ (
);

AND2X2 _18386_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_7296_)
);

FILL FILL_0__19462_ (
);

FILL FILL_0__19042_ (
);

FILL FILL182400x59280 (
);

FILL FILL_1__12976_ (
);

FILL FILL_1__12556_ (
);

FILL FILL_0__11969_ (
);

AND2X2 _11834_ (
    .A(_1734_),
    .B(_1733_),
    .Y(_1719_[7])
);

DFFSR _11414_ (
    .CLK(clk_bF$buf73),
    .D(_1455_[23]),
    .Q(\datapath_1.regfile_1.regOut[23] [23]),
    .R(rst_bF$buf39),
    .S(vdd)
);

FILL FILL_0__11129_ (
);

FILL FILL264480x39520 (
);

OR2X2 _12619_ (
    .A(_2183_),
    .B(_2181_),
    .Y(_2184_)
);

FILL FILL_1__17174_ (
);

OR2X2 _16872_ (
    .A(_5804_),
    .B(_5797_),
    .Y(_5805_)
);

FILL FILL_0__16167_ (
);

OR2X2 _16452_ (
    .A(_5389_),
    .B(_5390_),
    .Y(_5391_)
);

OR2X2 _16032_ (
    .A(_4977_),
    .B(_4974_),
    .Y(_4978_)
);

FILL FILL120840x74100 (
);

OR2X2 _8794_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .B(_200__bF$buf3),
    .Y(_188_)
);

FILL FILL_1__10202_ (
);

FILL FILL_1__18799_ (
);

FILL FILL279680x192660 (
);

FILL FILL207480x232180 (
);

OR2X2 _17657_ (
    .A(_6578_),
    .B(_6577_),
    .Y(_6579_)
);

AND2X2 _17237_ (
    .A(_4228__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_6164_)
);

NAND2X1 _12792_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2357_)
);

OR2X2 _12372_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_2013_)
);

FILL FILL_0__12087_ (
);

FILL FILL_0__18733_ (
);

FILL FILL107160x326040 (
);

FILL FILL_0__18313_ (
);

DFFSR _9999_ (
    .CLK(clk_bF$buf104),
    .D(_729_[27]),
    .Q(\datapath_1.regfile_1.regOut[12] [27]),
    .R(rst_bF$buf25),
    .S(vdd)
);

OR2X2 _9579_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_591_)
);

OR2X2 _9159_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_371_)
);

FILL FILL5320x54340 (
);

FILL FILL_0__8414_ (
);

FILL FILL503120x217360 (
);

FILL FILL_1__14299_ (
);

FILL FILL_0_BUFX2_insert790 (
);

FILL FILL_0_BUFX2_insert792 (
);

FILL FILL334400x212420 (
);

FILL FILL_0_BUFX2_insert793 (
);

OR2X2 _13997_ (
    .A(_3415_),
    .B(_3416_),
    .Y(_3417_)
);

FILL FILL_0_BUFX2_insert794 (
);

FILL FILL_0_BUFX2_insert795 (
);

OR2X2 _13577_ (
    .A(ALUOut[29]),
    .B(_3079__bF$buf1),
    .Y(_3073_)
);

NAND2X1 _13157_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(_2292_),
    .Y(_2708_)
);

FILL FILL_0_BUFX2_insert796 (
);

FILL FILL_0_BUFX2_insert797 (
);

FILL FILL_0_BUFX2_insert799 (
);

FILL FILL_0__19518_ (
);

FILL FILL345800x281580 (
);

FILL FILL211280x247000 (
);

FILL FILL28120x281580 (
);

FILL FILL161120x39520 (
);

FILL FILL_0__9619_ (
);

FILL FILL351120x128440 (
);

FILL FILL_1__16865_ (
);

FILL FILL342760x326040 (
);

FILL FILL_0__15438_ (
);

OR2X2 _15723_ (
    .A(_4672_),
    .B(_4673_),
    .Y(_4674_)
);

FILL FILL228760x350740 (
);

FILL FILL_0__15018_ (
);

OR2X2 _15303_ (
    .A(_4258_),
    .B(_4259_),
    .Y(_4260_)
);

FILL FILL_0__10573_ (
);

FILL FILL_0__10153_ (
);

AND2X2 _18195_ (
    .A(_6315__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_7108_)
);

FILL FILL168720x24700 (
);

FILL FILL414960x365560 (
);

FILL FILL9120x54340 (
);

FILL FILL_0__19271_ (
);

FILL FILL_1__12365_ (
);

OR2X2 _16928_ (
    .A(_5856_),
    .B(_5859_),
    .Y(_5860_)
);

AND2X2 _16508_ (
    .A(_4239__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_5446_)
);

FILL FILL_0__9792_ (
);

FILL FILL245480x266760 (
);

FILL FILL_0__11358_ (
);

OR2X2 _11643_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_1647_)
);

OR2X2 _11223_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_1427_)
);

FILL FILL_0__15191_ (
);

FILL FILL427880x177840 (
);

FILL FILL292600x54340 (
);

AND2X2 _12848_ (
    .A(_2412_),
    .B(_2410_),
    .Y(_2413_)
);

DFFSR _12428_ (
    .CLK(clk_bF$buf104),
    .D(_1983_[5]),
    .Q(\datapath_1.regfile_1.regOut[31] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

AND2X2 _12008_ (
    .A(_1830_),
    .B(_1829_),
    .Y(_1785_[22])
);

FILL FILL125400x340860 (
);

FILL FILL_0__13924_ (
);

FILL FILL_0__16396_ (
);

AND2X2 _16681_ (
    .A(_4217__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_5617_)
);

AND2X2 _16261_ (
    .A(_4195__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_5203_)
);

FILL FILL_1__15716_ (
);

FILL FILL_1__10011_ (
);

FILL FILL_1__18188_ (
);

OR2X2 _17886_ (
    .A(_6800_),
    .B(_6803_),
    .Y(_6804_)
);

OR2X2 _17466_ (
    .A(_6389_),
    .B(_6390_),
    .Y(_6391_)
);

OR2X2 _17046_ (
    .A(_5975_),
    .B(_5974_),
    .Y(_5976_)
);

DFFSR _12181_ (
    .CLK(clk_bF$buf76),
    .D(_1851_[16]),
    .Q(\datapath_1.regfile_1.regOut[29] [16]),
    .R(rst_bF$buf112),
    .S(vdd)
);

FILL FILL_0__18962_ (
);

FILL FILL_0__18542_ (
);

FILL FILL_0__18122_ (
);

FILL FILL87400x24700 (
);

OR2X2 _9388_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_530__bF$buf4),
    .Y(_484_)
);

FILL FILL478800x143260 (
);

FILL FILL169480x163020 (
);

FILL FILL_0__8643_ (
);

OR2X2 _10914_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_1261_)
);

FILL FILL_0__10209_ (
);

FILL FILL347320x251940 (
);

OR2X2 _13386_ (
    .A(_2397_),
    .B(_2376__bF$buf1),
    .Y(_2923_)
);

FILL FILL_0__19327_ (
);

FILL FILL_0__14462_ (
);

FILL FILL277400x256880 (
);

FILL FILL_0__14042_ (
);

FILL FILL_0__9428_ (
);

FILL FILL_0__9008_ (
);

FILL FILL427880x44460 (
);

FILL FILL241680x296400 (
);

FILL FILL64600x271700 (
);

OR2X2 _15952_ (
    .A(_4895_),
    .B(_4898_),
    .Y(_4899_)
);

FILL FILL_0__15667_ (
);

AND2X2 _15532_ (
    .A(_4225__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_4486_)
);

FILL FILL_0__15247_ (
);

AND2X2 _15112_ (
    .A(_4039_),
    .B(_4091_),
    .Y(_4092_)
);

FILL FILL23560x69160 (
);

FILL FILL55480x375440 (
);

FILL FILL_0__19080_ (
);

FILL FILL359480x286520 (
);

FILL FILL_1__17039_ (
);

FILL FILL118560x321100 (
);

FILL FILL235600x118560 (
);

AND2X2 _16737_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_5672_)
);

OR2X2 _16317_ (
    .A(_5257_),
    .B(_5256_),
    .Y(_5258_)
);

FILL FILL_0__11587_ (
);

OR2X2 _11872_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_1784__bF$buf4),
    .Y(_1760_)
);

OR2X2 _11452_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .B(_1586__bF$buf3),
    .Y(_1540_)
);

DFFSR _11032_ (
    .CLK(clk_bF$buf37),
    .D(_1257_[28]),
    .Q(\datapath_1.regfile_1.regOut[20] [28]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_0__17813_ (
);

FILL FILL499320x167960 (
);

OR2X2 _8659_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .B(_134__bF$buf3),
    .Y(_118_)
);

FILL FILL41040x202540 (
);

DFFSR _9600_ (
    .CLK(clk_bF$buf112),
    .D(_531_[15]),
    .Q(\datapath_1.regfile_1.regOut[9] [15]),
    .R(rst_bF$buf113),
    .S(vdd)
);

FILL FILL_1__13379_ (
);

XNOR2X1 _12657_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2222_)
);

OR2X2 _12237_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_1943_)
);

FILL FILL22040x360620 (
);

FILL FILL_1__14320_ (
);

FILL FILL457520x163020 (
);

FILL FILL44080x19760 (
);

FILL FILL129960x256880 (
);

FILL FILL_0__13313_ (
);

FILL FILL_0_BUFX2_insert1140 (
);

FILL FILL_0_BUFX2_insert1142 (
);

AND2X2 _16490_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_5429_)
);

AND2X2 _16070_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_5015_)
);

FILL FILL_0_BUFX2_insert1144 (
);

FILL FILL_0_BUFX2_insert1146 (
);

FILL FILL_0_BUFX2_insert1148 (
);

FILL FILL_0_BUFX2_insert1149 (
);

FILL FILL_1__15945_ (
);

AND2X2 _14803_ (
    .A(_3901_),
    .B(_3900_),
    .Y(_3870_[15])
);

AND2X2 _17695_ (
    .A(_6262__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_6616_)
);

INVX1 _17275_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_6201_)
);

FILL FILL_0__18771_ (
);

FILL FILL9120x365560 (
);

FILL FILL296400x370500 (
);

AND2X2 _9197_ (
    .A(_396_),
    .B(_395_),
    .Y(_333_[31])
);

FILL FILL_1__11865_ (
);

FILL FILL474240x266760 (
);

FILL FILL_0__8452_ (
);

FILL FILL_0__10858_ (
);

OR2X2 _10723_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .B(_1190__bF$buf1),
    .Y(_1174_)
);

FILL FILL_0__10018_ (
);

OR2X2 _10303_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .B(_992__bF$buf1),
    .Y(_954_)
);

AND2X2 _13195_ (
    .A(_2743_),
    .B(_2439_),
    .Y(_2744_)
);

OR2X2 _19421_ (
    .A(_8315_),
    .B(_8308_),
    .Y(_8316_)
);

FILL FILL_0__19136_ (
);

AND2X2 _19001_ (
    .A(_6272__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_7902_)
);

FILL FILL_0__14691_ (
);

FILL FILL_0__14271_ (
);

FILL FILL250800x311220 (
);

FILL FILL85880x69160 (
);

FILL FILL_0__9657_ (
);

DFFSR _11928_ (
    .CLK(clk_bF$buf34),
    .D(_1719_[21]),
    .Q(\datapath_1.regfile_1.regOut[27] [21]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_0__9237_ (
);

OR2X2 _11508_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_1577_)
);

FILL FILL374680x345800 (
);

FILL FILL248520x291460 (
);

FILL FILL422560x79040 (
);

FILL FILL_0__15896_ (
);

AND2X2 _15761_ (
    .A(_4187__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_4711_)
);

FILL FILL_0__15476_ (
);

AND2X2 _15341_ (
    .A(_4197__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_4298_)
);

FILL FILL_1__8613_ (
);

FILL FILL215080x79040 (
);

FILL FILL_1__17688_ (
);

FILL FILL_1__17268_ (
);

FILL FILL157320x34580 (
);

FILL FILL504640x167960 (
);

AND2X2 _16966_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_5897_)
);

AND2X2 _16546_ (
    .A(_4208__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_5484_)
);

AND2X2 _16126_ (
    .A(_4230__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_5070_)
);

OR2X2 _11681_ (
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .Y(_1717_)
);

AND2X2 _11261_ (
    .A(_1452_),
    .B(_1451_),
    .Y(_1389_[31])
);

FILL FILL_1__9818_ (
);

FILL FILL_0__17202_ (
);

AND2X2 _8888_ (
    .A(_230_),
    .B(_229_),
    .Y(_201_[14])
);

FILL FILL466640x29640 (
);

AND2X2 _8468_ (
    .A(_10_),
    .B(_9_),
    .Y(_3_[3])
);

FILL FILL297160x182780 (
);

NAND3X1 _12886_ (
    .A(_2273_),
    .B(_2269_),
    .C(_2270_),
    .Y(_2451_)
);

AND2X2 _12466_ (
    .A(_2051_),
    .B(_2058_),
    .Y(_2059_)
);

DFFSR _12046_ (
    .CLK(clk_bF$buf76),
    .D(_1785_[10]),
    .Q(\datapath_1.regfile_1.regOut[28] [10]),
    .R(rst_bF$buf112),
    .S(vdd)
);

FILL FILL_0__18827_ (
);

FILL FILL_0__18407_ (
);

FILL FILL_0__13962_ (
);

FILL FILL_0__13542_ (
);

FILL FILL_0__8928_ (
);

FILL FILL_0__8508_ (
);

FILL FILL470440x296400 (
);

FILL FILL159600x242060 (
);

FILL FILL304760x9880 (
);

FILL FILL_1__15334_ (
);

FILL FILL115520x64220 (
);

DFFSR _14612_ (
    .CLK(clk_bF$buf15),
    .D(_3738_[18]),
    .Q(\datapath_1.PCJump [20]),
    .R(rst_bF$buf31),
    .S(vdd)
);

FILL FILL_0__14327_ (
);

FILL FILL12160x103740 (
);

AND2X2 _17084_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_6013_)
);

FILL FILL_0__18580_ (
);

FILL FILL_0__18160_ (
);

FILL FILL_1__11254_ (
);

OR2X2 _15817_ (
    .A(_4765_),
    .B(_4758_),
    .Y(_4766_)
);

FILL FILL123880x148200 (
);

FILL FILL192280x34580 (
);

FILL FILL_0__8681_ (
);

AND2X2 _10952_ (
    .A(_1286_),
    .B(_1285_),
    .Y(_1257_[14])
);

FILL FILL_0__10667_ (
);

AND2X2 _10532_ (
    .A(_1066_),
    .B(_1065_),
    .Y(_1059_[3])
);

DFFSR _10112_ (
    .CLK(clk_bF$buf57),
    .D(_795_[11]),
    .Q(\datapath_1.regfile_1.regOut[13] [11]),
    .R(rst_bF$buf39),
    .S(vdd)
);

FILL FILL246240x340860 (
);

FILL FILL76000x34580 (
);

OR2X2 _18289_ (
    .A(_7199_),
    .B(_7200_),
    .Y(_7201_)
);

FILL FILL77520x242060 (
);

AND2X2 _19230_ (
    .A(_8127_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.rd1 [28])
);

FILL FILL484880x79040 (
);

FILL FILL349600x365560 (
);

FILL FILL244720x187720 (
);

OR2X2 _11737_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .B(_1718__bF$buf2),
    .Y(_1690_)
);

FILL FILL_0__9046_ (
);

OR2X2 _11317_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .B(_1520__bF$buf2),
    .Y(_1470_)
);

FILL FILL_1__13820_ (
);

FILL FILL446880x316160 (
);

FILL FILL_0__12813_ (
);

FILL FILL_1__16292_ (
);

FILL FILL436240x276640 (
);

FILL FILL230280x49400 (
);

OR2X2 _15990_ (
    .A(_4933_),
    .B(_4936_),
    .Y(_4937_)
);

FILL FILL_0__15285_ (
);

AND2X2 _15570_ (
    .A(_4208__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_4523_)
);

NOR2X1 _15150_ (
    .A(_4080_),
    .B(_4042_),
    .Y(\datapath_1.regfile_1.regEn [24])
);

FILL FILL_1__8422_ (
);

FILL FILL197600x276640 (
);

OR2X2 _16775_ (
    .A(_5707_),
    .B(_5708_),
    .Y(_5709_)
);

OR2X2 _16355_ (
    .A(_5294_),
    .B(_5295_),
    .Y(_5296_)
);

OR2X2 _11490_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_1565_)
);

OR2X2 _11070_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_1345_)
);

FILL FILL_1__9627_ (
);

FILL FILL_0__17851_ (
);

FILL FILL_0__17431_ (
);

FILL FILL257640x49400 (
);

DFFSR _8697_ (
    .CLK(clk_bF$buf90),
    .D(_69_[15]),
    .Q(\datapath_1.regfile_1.regOut[2] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL_1__10945_ (
);

FILL FILL180880x345800 (
);

BUFX2 BUFX2_insert390 (
    .A(_6259_),
    .Y(_6259__bF$buf0)
);

BUFX2 BUFX2_insert391 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf4 )
);

BUFX2 BUFX2_insert392 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf3 )
);

BUFX2 BUFX2_insert393 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf2 )
);

BUFX2 BUFX2_insert394 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf1 )
);

BUFX2 BUFX2_insert395 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf0 )
);

BUFX2 BUFX2_insert396 (
    .A(_6297_),
    .Y(_6297__bF$buf4)
);

BUFX2 BUFX2_insert397 (
    .A(_6297_),
    .Y(_6297__bF$buf3)
);

BUFX2 BUFX2_insert398 (
    .A(_6297_),
    .Y(_6297__bF$buf2)
);

INVX1 _12695_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .Y(_2260_)
);

BUFX2 BUFX2_insert399 (
    .A(_6297_),
    .Y(_6297__bF$buf1)
);

AND2X2 _12275_ (
    .A(_1968_),
    .B(_1967_),
    .Y(_1917_[25])
);

FILL FILL_0__18636_ (
);

AND2X2 _18921_ (
    .A(_6244__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_7823_)
);

AND2X2 _18501_ (
    .A(_6232__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_7410_)
);

FILL FILL417240x222300 (
);

FILL FILL_0__13771_ (
);

FILL FILL91960x93860 (
);

FILL FILL_0__8737_ (
);

FILL FILL411160x375440 (
);

FILL FILL38000x64220 (
);

FILL FILL_0__14976_ (
);

OR2X2 _14841_ (
    .A(\datapath_1.rd2 [28]),
    .B(_3935__bF$buf4),
    .Y(_3927_)
);

FILL FILL_0__14136_ (
);

OR2X2 _14421_ (
    .A(memoryOutData[17]),
    .B(_3737__bF$buf3),
    .Y(_3707_)
);

OR2X2 _14001_ (
    .A(_3420_),
    .B(_3417_),
    .Y(\datapath_1.alu_1.ALUInB [11])
);

FILL FILL233320x345800 (
);

FILL FILL_1__11063_ (
);

FILL FILL73720x138320 (
);

AND2X2 _15626_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_4578_)
);

FILL FILL198360x14820 (
);

OR2X2 _15206_ (
    .A(_4149_),
    .B(_4163_),
    .Y(_4164_)
);

FILL FILL_0__8490_ (
);

FILL FILL_0__10476_ (
);

DFFSR _10761_ (
    .CLK(clk_bF$buf89),
    .D(_1125_[15]),
    .Q(\datapath_1.regfile_1.regOut[18] [15]),
    .R(rst_bF$buf83),
    .S(vdd)
);

OR2X2 _10341_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_979_)
);

FILL FILL_0__10056_ (
);

OR2X2 _18098_ (
    .A(_7012_),
    .B(_7009_),
    .Y(_7013_)
);

FILL FILL_0__16702_ (
);

FILL FILL477280x182780 (
);

FILL FILL_0__19174_ (
);

FILL FILL_1__12268_ (
);

FILL FILL_0__9695_ (
);

AND2X2 _11966_ (
    .A(_1802_),
    .B(_1801_),
    .Y(_1785_[8])
);

DFFSR _11546_ (
    .CLK(clk_bF$buf86),
    .D(_1521_[26]),
    .Q(\datapath_1.regfile_1.regOut[24] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

FILL FILL90440x375440 (
);

AND2X2 _11126_ (
    .A(_1382_),
    .B(_1381_),
    .Y(_1323_[29])
);

FILL FILL_0__17907_ (
);

FILL FILL_0__12202_ (
);

FILL FILL_0__15094_ (
);

FILL FILL348840x133380 (
);

FILL FILL234080x291460 (
);

FILL FILL_0__13827_ (
);

FILL FILL_0__13407_ (
);

OR2X2 _16584_ (
    .A(_5520_),
    .B(_5517_),
    .Y(_5521_)
);

AND2X2 _16164_ (
    .A(_4217__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_5108_)
);

FILL FILL_1__9016_ (
);

FILL FILL_0__17660_ (
);

FILL FILL284240x306280 (
);

FILL FILL_0__17240_ (
);

FILL FILL_1__10334_ (
);

FILL FILL270560x330980 (
);

FILL FILL238640x172900 (
);

AND2X2 _17789_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_6709_)
);

INVX1 _17369_ (
    .A(_6257_),
    .Y(_6295_)
);

FILL FILL_1__19452_ (
);

OR2X2 _12084_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_1861_)
);

FILL FILL288040x227240 (
);

OR2X2 _18730_ (
    .A(_7633_),
    .B(_7634_),
    .Y(_7635_)
);

AND2X2 _18310_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_7222_)
);

FILL FILL_0__18025_ (
);

FILL FILL_0__13580_ (
);

FILL FILL_0__13160_ (
);

FILL FILL_1__11959_ (
);

AND2X2 _10817_ (
    .A(_1216_),
    .B(_1215_),
    .Y(_1191_[12])
);

FILL FILL122360x158080 (
);

AND2X2 _13289_ (
    .A(_2791_),
    .B(_2831_),
    .Y(_2832_)
);

OR2X2 _19515_ (
    .A(gnd),
    .B(_8385__bF$buf0),
    .Y(_8379_)
);

FILL FILL_0__14785_ (
);

AND2X2 _14650_ (
    .A(_3819_),
    .B(_3818_),
    .Y(_3804_[7])
);

OR2X2 _14230_ (
    .A(MemToReg_bF$buf4),
    .B(ALUOut[29]),
    .Y(_3598_)
);

FILL FILL23560x242060 (
);

FILL FILL503120x34580 (
);

FILL FILL327560x153140 (
);

FILL FILL_1__16157_ (
);

FILL FILL101840x83980 (
);

FILL FILL14440x217360 (
);

OR2X2 _15855_ (
    .A(_4800_),
    .B(_4803_),
    .Y(_4804_)
);

AND2X2 _15435_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_4390_)
);

NOR3X1 _15015_ (
    .A(_4003_),
    .B(\datapath_1.a3 [1]),
    .C(_4002_),
    .Y(_4004_)
);

FILL FILL413440x69160 (
);

FILL FILL266000x281580 (
);

OR2X2 _10990_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .B(_1322__bF$buf4),
    .Y(_1312_)
);

FILL FILL_0__10285_ (
);

OR2X2 _10570_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .B(_1124__bF$buf1),
    .Y(_1092_)
);

OR2X2 _10150_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .B(_926__bF$buf3),
    .Y(_872_)
);

FILL FILL_0__16931_ (
);

FILL FILL380760x242060 (
);

OR2X2 _11775_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_1715_)
);

OR2X2 _11355_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_1495_)
);

FILL FILL98040x88920 (
);

FILL FILL55480x4940 (
);

FILL FILL_0__17716_ (
);

FILL FILL13680x14820 (
);

AND2X2 _9923_ (
    .A(_760_),
    .B(_759_),
    .Y(_729_[15])
);

AND2X2 _9503_ (
    .A(_540_),
    .B(_539_),
    .Y(_531_[4])
);

FILL FILL147440x197600 (
);

FILL FILL380760x108680 (
);

FILL FILL417240x69160 (
);

FILL FILL253080x271700 (
);

AND2X2 _13921_ (
    .A(ALUSrcB[0]),
    .B(ALUSrcB[1]),
    .Y(_3352_)
);

FILL FILL_0__13636_ (
);

OR2X2 _13501_ (
    .A(IorD_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [4]),
    .Y(_3022_)
);

FILL FILL80560x118560 (
);

OR2X2 _16393_ (
    .A(_5325_),
    .B(_5332_),
    .Y(_5333_)
);

FILL FILL_1__10143_ (
);

OR2X2 _14706_ (
    .A(\datapath_1.rd1 [26]),
    .B(_3869__bF$buf0),
    .Y(_3857_)
);

BUFX2 BUFX2_insert770 (
    .A(_6229_),
    .Y(_6229__bF$buf2)
);

BUFX2 BUFX2_insert771 (
    .A(_6229_),
    .Y(_6229__bF$buf1)
);

BUFX2 BUFX2_insert772 (
    .A(_6229_),
    .Y(_6229__bF$buf0)
);

BUFX2 BUFX2_insert773 (
    .A(_1784_),
    .Y(_1784__bF$buf4)
);

FILL FILL84360x360620 (
);

BUFX2 BUFX2_insert774 (
    .A(_1784_),
    .Y(_1784__bF$buf3)
);

AND2X2 _17598_ (
    .A(_6236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_6521_)
);

BUFX2 BUFX2_insert775 (
    .A(_1784_),
    .Y(_1784__bF$buf2)
);

BUFX2 BUFX2_insert776 (
    .A(_1784_),
    .Y(_1784__bF$buf1)
);

AND2X2 _17178_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_6106_)
);

BUFX2 BUFX2_insert777 (
    .A(_1784_),
    .Y(_1784__bF$buf0)
);

BUFX2 BUFX2_insert778 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf4 )
);

BUFX2 BUFX2_insert779 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf3 )
);

FILL FILL65360x197600 (
);

FILL FILL37240x29640 (
);

FILL FILL_0__18674_ (
);

FILL FILL_0__18254_ (
);

FILL FILL160360x301340 (
);

FILL FILL_0__8775_ (
);

FILL FILL10640x247000 (
);

DFFSR _10626_ (
    .CLK(clk_bF$buf75),
    .D(_1059_[9]),
    .Q(\datapath_1.regfile_1.regOut[17] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

OR2X2 _10206_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_909_)
);

AND2X2 _13098_ (
    .A(_2652_),
    .B(_2639_),
    .Y(_2653_)
);

FILL FILL_0__19039_ (
);

OR2X2 _19324_ (
    .A(_8212_),
    .B(_8219_),
    .Y(_8220_)
);

FILL FILL_0__12907_ (
);

FILL FILL_1__16386_ (
);

FILL FILL295640x301340 (
);

FILL FILL_0__15379_ (
);

AND2X2 _15664_ (
    .A(_4208__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_4616_)
);

AND2X2 _15244_ (
    .A(_4171_),
    .B(_4165_),
    .Y(_4202_)
);

FILL FILL_0__10094_ (
);

FILL FILL481840x316160 (
);

FILL FILL_0__16320_ (
);

AND2X2 _16869_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_5802_)
);

OR2X2 _16449_ (
    .A(_5387_),
    .B(_5384_),
    .Y(_5388_)
);

AND2X2 _16029_ (
    .A(_4187__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_4975_)
);

FILL FILL82080x222300 (
);

FILL FILL228760x24700 (
);

OR2X2 _11584_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .B(_1652__bF$buf4),
    .Y(_1608_)
);

DFFSR _11164_ (
    .CLK(clk_bF$buf111),
    .D(_1323_[31]),
    .Q(\datapath_1.regfile_1.regOut[21] [31]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL479560x69160 (
);

FILL FILL_0__17945_ (
);

FILL FILL_0__17525_ (
);

AND2X2 _17810_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_6729_)
);

FILL FILL_0__17105_ (
);

FILL FILL_0__12660_ (
);

FILL FILL_0__12240_ (
);

FILL FILL451440x9880 (
);

FILL FILL297920x0 (
);

FILL FILL432440x39520 (
);

DFFSR _9732_ (
    .CLK(clk_bF$buf103),
    .D(_597_[18]),
    .Q(\datapath_1.regfile_1.regOut[10] [18]),
    .R(rst_bF$buf45),
    .S(vdd)
);

OR2X2 _9312_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_453_)
);

NAND2X1 _12789_ (
    .A(_2351_),
    .B(_2352_),
    .Y(_2354_)
);

OR2X2 _12369_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_2011_)
);

FILL FILL_1__19317_ (
);

FILL FILL503120x330980 (
);

FILL FILL_1__14452_ (
);

FILL FILL_0__13865_ (
);

FILL FILL_0__13445_ (
);

OR2X2 _13730_ (
    .A(_3205_),
    .B(_3202_),
    .Y(\datapath_1.mux_pcsrc.dout [19])
);

FILL FILL_0__13025_ (
);

AND2X2 _13310_ (
    .A(_2850_),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2851_)
);

FILL FILL434720x4940 (
);

FILL FILL_1__9054_ (
);

FILL FILL446120x281580 (
);

FILL FILL412680x113620 (
);

AND2X2 _14935_ (
    .A(_3969_),
    .B(_3968_),
    .Y(_3936_[16])
);

AND2X2 _14515_ (
    .A(_3749_),
    .B(_3748_),
    .Y(_3738_[5])
);

FILL FILL453720x4940 (
);

FILL FILL_1__19070_ (
);

FILL FILL181640x44460 (
);

FILL FILL_1__11997_ (
);

FILL FILL346560x360620 (
);

OR2X2 _10855_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .B(_1256__bF$buf2),
    .Y(_1242_)
);

OR2X2 _10435_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .B(_1058__bF$buf3),
    .Y(_1022_)
);

OR2X2 _10015_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .B(_860__bF$buf1),
    .Y(_802_)
);

FILL FILL86640x83980 (
);

FILL FILL_0__19268_ (
);

DFFSR _19553_ (
    .CLK(clk_bF$buf33),
    .D(_8320_[30]),
    .Q(\datapath_1.regfile_1.regOut[0] [30]),
    .R(rst_bF$buf88),
    .S(vdd)
);

OR2X2 _19133_ (
    .A(_8030_),
    .B(_8031_),
    .Y(_8032_)
);

FILL FILL_0__9789_ (
);

FILL FILL_0__9369_ (
);

FILL FILL300960x301340 (
);

FILL FILL_1__13303_ (
);

AND2X2 _15893_ (
    .A(_4223__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_4841_)
);

AND2X2 _15473_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_4428_)
);

NAND2X1 _15053_ (
    .A(\datapath_1.a3 [4]),
    .B(RegWrite),
    .Y(_4042_)
);

FILL FILL_1__8745_ (
);

FILL FILL_1__14508_ (
);

FILL FILL494760x39520 (
);

FILL FILL383800x133380 (
);

OR2X2 _16678_ (
    .A(_5613_),
    .B(_5612_),
    .Y(_5614_)
);

AND2X2 _16258_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_5200_)
);

DFFSR _11393_ (
    .CLK(clk_bF$buf17),
    .D(_1455_[2]),
    .Q(\datapath_1.regfile_1.regOut[23] [2]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL287280x39520 (
);

FILL FILL_0__17754_ (
);

FILL FILL302480x296400 (
);

OR2X2 _9961_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .B(_794__bF$buf1),
    .Y(_786_)
);

OR2X2 _9541_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_596__bF$buf4),
    .Y(_566_)
);

OR2X2 _9121_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .B(_398__bF$buf3),
    .Y(_346_)
);

NAND2X1 _12598_ (
    .A(\datapath_1.alu_1.ALUInA [30]),
    .B(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2163_)
);

DFFSR _12178_ (
    .CLK(clk_bF$buf4),
    .D(_1851_[13]),
    .Q(\datapath_1.regfile_1.regOut[29] [13]),
    .R(rst_bF$buf70),
    .S(vdd)
);

FILL FILL_1__14261_ (
);

OR2X2 _18824_ (
    .A(_7727_),
    .B(_7726_),
    .Y(_7728_)
);

FILL FILL_0__18539_ (
);

FILL FILL_0__18119_ (
);

FILL FILL_0_BUFX2_insert411 (
);

OR2X2 _18404_ (
    .A(_7313_),
    .B(_7312_),
    .Y(_7314_)
);

FILL FILL_0_BUFX2_insert413 (
);

FILL FILL_0_BUFX2_insert414 (
);

FILL FILL_0__13254_ (
);

FILL FILL_0_BUFX2_insert415 (
);

FILL FILL_0_BUFX2_insert416 (
);

FILL FILL481840x93860 (
);

FILL FILL_0_BUFX2_insert417 (
);

FILL FILL_0_BUFX2_insert419 (
);

FILL FILL370880x123500 (
);

FILL FILL_1__15886_ (
);

FILL FILL209760x232180 (
);

DFFSR _14744_ (
    .CLK(clk_bF$buf38),
    .D(_3804_[21]),
    .Q(\datapath_1.a [21]),
    .R(rst_bF$buf70),
    .S(vdd)
);

FILL FILL_0__14459_ (
);

OR2X2 _14324_ (
    .A(vdd),
    .B(ALUOut[28]),
    .Y(_3662_)
);

FILL FILL437760x296400 (
);

FILL FILL_0__15820_ (
);

FILL FILL_0__15400_ (
);

FILL FILL287280x360620 (
);

FILL FILL_0__18292_ (
);

FILL FILL488680x113620 (
);

FILL FILL316920x19760 (
);

FILL FILL505400x217360 (
);

FILL FILL_1__11386_ (
);

AND2X2 _15949_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_4896_)
);

AND2X2 _15529_ (
    .A(_4234__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_4483_)
);

AND2X2 _15109_ (
    .A(_4029_),
    .B(_4089_),
    .Y(\datapath_1.regfile_1.regEn [9])
);

FILL FILL_0__8393_ (
);

FILL FILL_0__10799_ (
);

AND2X2 _10664_ (
    .A(_1134_),
    .B(_1133_),
    .Y(_1125_[4])
);

DFFSR _10244_ (
    .CLK(clk_bF$buf1),
    .D(_861_[14]),
    .Q(\datapath_1.regfile_1.regOut[14] [14]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL164160x24700 (
);

FILL FILL109440x19760 (
);

FILL FILL250040x103740 (
);

FILL FILL_0__19497_ (
);

FILL FILL278160x93860 (
);

AND2X2 _19362_ (
    .A(_6328__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_8257_)
);

FILL FILL_0__19077_ (
);

FILL FILL180120x108680 (
);

DFFSR _8812_ (
    .CLK(clk_bF$buf1),
    .D(_135_[1]),
    .Q(\datapath_1.regfile_1.regOut[3] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

FILL FILL_0__9178_ (
);

OR2X2 _11869_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .B(_1784__bF$buf2),
    .Y(_1758_)
);

OR2X2 _11449_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .B(_1586__bF$buf3),
    .Y(_1538_)
);

DFFSR _11029_ (
    .CLK(clk_bF$buf41),
    .D(_1257_[25]),
    .Q(\datapath_1.regfile_1.regOut[20] [25]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL_1__13952_ (
);

FILL FILL_0__12945_ (
);

OR2X2 _12810_ (
    .A(ALUControl[1]),
    .B(ALUControl[0]),
    .Y(_2375_)
);

FILL FILL_0__12525_ (
);

FILL FILL_0__12105_ (
);

AND2X2 _15282_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_4240_)
);

FILL FILL256880x291460 (
);

FILL FILL357200x370500 (
);

FILL FILL348840x247000 (
);

OR2X2 _16487_ (
    .A(_5425_),
    .B(_5422_),
    .Y(_5426_)
);

AND2X2 _16067_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_5012_)
);

FILL FILL_1__18570_ (
);

FILL FILL_1__18150_ (
);

FILL FILL_1__9759_ (
);

FILL FILL_0__17143_ (
);

AND2X2 _9770_ (
    .A(_678_),
    .B(_677_),
    .Y(_663_[7])
);

DFFSR _9350_ (
    .CLK(clk_bF$buf87),
    .D(_399_[23]),
    .Q(\datapath_1.regfile_1.regOut[7] [23]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL11400x321100 (
);

FILL FILL_0__18768_ (
);

OR2X2 _18633_ (
    .A(_7539_),
    .B(_7536_),
    .Y(_7540_)
);

FILL FILL_0__18348_ (
);

OR2X2 _18213_ (
    .A(_7125_),
    .B(_7124_),
    .Y(_7126_)
);

FILL FILL_0__13483_ (
);

FILL FILL_0__8869_ (
);

FILL FILL_0__8449_ (
);

FILL FILL_1__12803_ (
);

FILL FILL97280x148200 (
);

FILL FILL_0__9810_ (
);

FILL FILL_1__15275_ (
);

AND2X2 _19418_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_8313_)
);

OR2X2 _14973_ (
    .A(\datapath_1.mux_pcsrc.dout [29]),
    .B(_4001__bF$buf3),
    .Y(_3995_)
);

FILL FILL_0__14268_ (
);

OR2X2 _14553_ (
    .A(memoryOutData[18]),
    .B(_3803__bF$buf4),
    .Y(_3775_)
);

OR2X2 _14133_ (
    .A(_3533_),
    .B(_3532_),
    .Y(_3534_)
);

FILL FILL154280x247000 (
);

FILL FILL_1__11195_ (
);

FILL FILL349600x251940 (
);

AND2X2 _15758_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_4708_)
);

AND2X2 _15338_ (
    .A(_4239__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_4295_)
);

DFFSR _10893_ (
    .CLK(clk_bF$buf37),
    .D(_1191_[18]),
    .Q(\datapath_1.regfile_1.regOut[19] [18]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL_0__10188_ (
);

OR2X2 _10473_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_1047_)
);

OR2X2 _10053_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_827_)
);

FILL FILL_0__16834_ (
);

FILL FILL_0__16414_ (
);

FILL FILL226480x286520 (
);

FILL FILL375440x192660 (
);

OR2X2 _19171_ (
    .A(_8068_),
    .B(_8067_),
    .Y(_8069_)
);

FILL FILL467400x148200 (
);

AND2X2 _8621_ (
    .A(_92_),
    .B(_91_),
    .Y(_69_[11])
);

FILL FILL453720x172900 (
);

DFFSR _11678_ (
    .CLK(clk_bF$buf107),
    .D(_1587_[29]),
    .Q(\datapath_1.regfile_1.regOut[25] [29]),
    .R(rst_bF$buf37),
    .S(vdd)
);

AND2X2 _11258_ (
    .A(_1450_),
    .B(_1449_),
    .Y(_1389_[30])
);

FILL FILL_0__17619_ (
);

AND2X2 _17904_ (
    .A(_6221__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_6822_)
);

FILL FILL_0__12754_ (
);

FILL FILL_0__12334_ (
);

NAND3X1 _15091_ (
    .A(_4020_),
    .B(_4054_),
    .C(_4017_),
    .Y(_4075_)
);

OR2X2 _9826_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .B(_728__bF$buf0),
    .Y(_716_)
);

OR2X2 _9406_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .B(_530__bF$buf2),
    .Y(_496_)
);

FILL FILL438520x232180 (
);

FILL FILL_1__14126_ (
);

FILL FILL_0__13959_ (
);

AND2X2 _13824_ (
    .A(_3282_),
    .B(_3281_),
    .Y(\datapath_1.alu_1.ALUInA [2])
);

FILL FILL_0__13119_ (
);

OR2X2 _13404_ (
    .A(_2939_),
    .B(_2376__bF$buf1),
    .Y(_2940_)
);

FILL FILL133760x316160 (
);

FILL FILL82840x59280 (
);

OR2X2 _16296_ (
    .A(_5230_),
    .B(_5237_),
    .Y(_5238_)
);

FILL FILL_0__14900_ (
);

FILL FILL_1__9148_ (
);

FILL FILL_0__17792_ (
);

FILL FILL_0__17372_ (
);

FILL FILL140600x286520 (
);

DFFSR _14609_ (
    .CLK(clk_bF$buf58),
    .D(_3738_[15]),
    .Q(\datapath_1.PCJump [17]),
    .R(rst_bF$buf15),
    .S(vdd)
);

FILL FILL24320x360620 (
);

FILL FILL_0__10820_ (
);

FILL FILL317680x49400 (
);

FILL FILL_0__18997_ (
);

AND2X2 _18862_ (
    .A(_6293__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_7765_)
);

FILL FILL_0__18157_ (
);

AND2X2 _18442_ (
    .A(_6287__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_7352_)
);

FILL FILL237880x330980 (
);

FILL FILL319960x148200 (
);

OR2X2 _18022_ (
    .A(_6937_),
    .B(_6934_),
    .Y(_6938_)
);

AND2X2 _10949_ (
    .A(_1284_),
    .B(_1283_),
    .Y(_1257_[13])
);

AND2X2 _10529_ (
    .A(_1064_),
    .B(_1063_),
    .Y(_1059_[2])
);

DFFSR _10109_ (
    .CLK(clk_bF$buf61),
    .D(_795_[8]),
    .Q(\datapath_1.regfile_1.regOut[13] [8]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL355680x227240 (
);

FILL FILL_0__11605_ (
);

FILL FILL463600x19760 (
);

OR2X2 _19227_ (
    .A(_8108_),
    .B(_8124_),
    .Y(_8125_)
);

AND2X2 _14782_ (
    .A(_3887_),
    .B(_3886_),
    .Y(_3870_[8])
);

FILL FILL_0__14077_ (
);

DFFSR _14362_ (
    .CLK(clk_bF$buf41),
    .D(_3606_[26]),
    .Q(ALUOut[26]),
    .R(rst_bF$buf63),
    .S(vdd)
);

FILL FILL381520x360620 (
);

FILL FILL441560x79040 (
);

FILL FILL164160x9880 (
);

AND2X2 _15987_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_4934_)
);

OR2X2 _15567_ (
    .A(_4519_),
    .B(_4518_),
    .Y(_4520_)
);

AND2X2 _15147_ (
    .A(_4110_),
    .B(_4113_),
    .Y(_4114_)
);

OR2X2 _10282_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_992__bF$buf4),
    .Y(_940_)
);

FILL FILL_0__16643_ (
);

FILL FILL499320x350740 (
);

FILL FILL421800x316160 (
);

FILL FILL_0__16223_ (
);

FILL FILL322240x212420 (
);

OR2X2 _8850_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_205_)
);

BUFX2 _8430_ (
    .A(_2_[6]),
    .Y(memoryWriteData[6])
);

OR2X2 _11487_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_1563_)
);

FILL FILL_1__18435_ (
);

OR2X2 _11067_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_1343_)
);

FILL FILL_1__18015_ (
);

FILL FILL376960x345800 (
);

FILL FILL421800x49400 (
);

FILL FILL59280x345800 (
);

FILL FILL445360x79040 (
);

AND2X2 _17713_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_6634_)
);

FILL FILL462080x29640 (
);

FILL FILL_0__17008_ (
);

FILL FILL_0__12983_ (
);

FILL FILL166440x4940 (
);

AND2X2 _9635_ (
    .A(_608_),
    .B(_607_),
    .Y(_597_[5])
);

DFFSR _9215_ (
    .CLK(clk_bF$buf6),
    .D(_333_[17]),
    .Q(\datapath_1.regfile_1.regOut[6] [17]),
    .R(rst_bF$buf31),
    .S(vdd)
);

OR2X2 _18918_ (
    .A(_7818_),
    .B(_7819_),
    .Y(_7820_)
);

FILL FILL_0__13348_ (
);

AND2X2 _13633_ (
    .A(_3081__bF$buf2),
    .B(ALUOut[6]),
    .Y(_3122_)
);

AND2X2 _13213_ (
    .A(_2760_),
    .B(_2547_),
    .Y(_2761_)
);

FILL FILL_1__10695_ (
);

FILL FILL299440x182780 (
);

OR2X2 _14838_ (
    .A(\datapath_1.rd2 [27]),
    .B(_3935__bF$buf2),
    .Y(_3925_)
);

OR2X2 _14418_ (
    .A(memoryOutData[16]),
    .B(_3737__bF$buf3),
    .Y(_3705_)
);

FILL FILL_0__15914_ (
);

FILL FILL446880x88920 (
);

AND2X2 _18671_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_7577_)
);

FILL FILL_0__18386_ (
);

OR2X2 _18251_ (
    .A(_7156_),
    .B(_7163_),
    .Y(_7164_)
);

FILL FILL386080x44460 (
);

FILL FILL_0__8487_ (
);

DFFSR _10758_ (
    .CLK(clk_bF$buf103),
    .D(_1125_[12]),
    .Q(\datapath_1.regfile_1.regOut[18] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

OR2X2 _10338_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_977_)
);

FILL FILL500840x108680 (
);

AND2X2 _19456_ (
    .A(_8339_),
    .B(_8338_),
    .Y(_8320_[9])
);

AND2X2 _19036_ (
    .A(_6300__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_7936_)
);

OR2X2 _14591_ (
    .A(IRWrite_bF$buf2),
    .B(\control_1.op [5]),
    .Y(_3800_)
);

OR2X2 _14171_ (
    .A(\datapath_1.Data [9]),
    .B(_3605__bF$buf0),
    .Y(_3559_)
);

AND2X2 _8906_ (
    .A(_242_),
    .B(_241_),
    .Y(_201_[20])
);

FILL FILL452200x182780 (
);

FILL FILL_1__13626_ (
);

OR2X2 _12904_ (
    .A(_2466_),
    .B(_2468_),
    .Y(_2469_)
);

FILL FILL_0__12619_ (
);

FILL FILL504640x350740 (
);

FILL FILL_1_BUFX2_insert345 (
);

FILL FILL_1_BUFX2_insert347 (
);

FILL FILL_1_BUFX2_insert349 (
);

AND2X2 _15796_ (
    .A(_4177__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_4746_)
);

OR2X2 _15376_ (
    .A(_4328_),
    .B(_4331_),
    .Y(_4332_)
);

AND2X2 _10091_ (
    .A(_852_),
    .B(_851_),
    .Y(_795_[28])
);

FILL FILL_1__8648_ (
);

FILL FILL_0__16872_ (
);

FILL FILL_1__18664_ (
);

OR2X2 _11296_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(_1520__bF$buf0),
    .Y(_1456_)
);

AND2X2 _17942_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_6859_)
);

FILL FILL_0__17657_ (
);

FILL FILL_0__17237_ (
);

AND2X2 _17522_ (
    .A(_6287__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_6446_)
);

AND2X2 _17102_ (
    .A(_4175__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_6031_)
);

DFFSR _9864_ (
    .CLK(clk_bF$buf28),
    .D(_663_[21]),
    .Q(\datapath_1.regfile_1.regOut[11] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

OR2X2 _9444_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_521_)
);

OR2X2 _9024_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_301_)
);

FILL FILL_1__14584_ (
);

FILL FILL118560x59280 (
);

AND2X2 _18727_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_7632_)
);

OR2X2 _18307_ (
    .A(_7217_),
    .B(_7218_),
    .Y(_7219_)
);

FILL FILL_0__13997_ (
);

OR2X2 _13862_ (
    .A(\datapath_1.a [15]),
    .B(_3342__bF$buf0),
    .Y(_3308_)
);

FILL FILL_0__13577_ (
);

AND2X2 _13442_ (
    .A(_2684_),
    .B(_2653_),
    .Y(_2975_)
);

OAI21X1 _13022_ (
    .A(_2286_),
    .B(_2259_),
    .C(_2316_),
    .Y(_2581_)
);

FILL FILL348080x74100 (
);

FILL FILL_1__15369_ (
);

FILL FILL_1__10084_ (
);

FILL FILL502360x212420 (
);

AND2X2 _14647_ (
    .A(_3817_),
    .B(_3816_),
    .Y(_3804_[6])
);

FILL FILL240920x128440 (
);

FILL FILL454480x0 (
);

OR2X2 _14227_ (
    .A(MemToReg_bF$buf1),
    .B(ALUOut[28]),
    .Y(_3596_)
);

FILL FILL_0__15303_ (
);

FILL FILL329840x59280 (
);

FILL FILL_0__18195_ (
);

OR2X2 _18480_ (
    .A(_7388_),
    .B(_7374_),
    .Y(_7389_)
);

AND2X2 _18060_ (
    .A(_6975_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd1 [10])
);

FILL FILL208240x197600 (
);

FILL FILL413440x375440 (
);

OR2X2 _10987_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .B(_1322__bF$buf4),
    .Y(_1310_)
);

FILL FILL_1__17515_ (
);

OR2X2 _10567_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_1124__bF$buf4),
    .Y(_1090_)
);

OR2X2 _10147_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .B(_926__bF$buf1),
    .Y(_870_)
);

FILL FILL_0__16508_ (
);

FILL FILL_0__11223_ (
);

AND2X2 _19265_ (
    .A(_6312__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_8162_)
);

INVX2 _8715_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .Y(_200_)
);

FILL FILL202920x44460 (
);

FILL FILL_0__12848_ (
);

NAND2X1 _12713_ (
    .A(\datapath_1.alu_1.ALUInA [19]),
    .B(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2278_)
);

FILL FILL_0__12008_ (
);

AND2X2 _15185_ (
    .A(_4142__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_4143_)
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_1_BUFX2_insert19 (
);

FILL FILL_1__8457_ (
);

FILL FILL_0__16261_ (
);

FILL FILL342000x153140 (
);

FILL FILL379240x276640 (
);

OR2X2 _13918_ (
    .A(_3345_),
    .B(_3348_),
    .Y(_3349_)
);

FILL FILL396720x286520 (
);

FILL FILL79040x286520 (
);

FILL FILL206720x44460 (
);

FILL FILL_0__17886_ (
);

FILL FILL_0__17466_ (
);

OR2X2 _17751_ (
    .A(_6662_),
    .B(_6670_),
    .Y(_6671_)
);

OR2X2 _17331_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_6257_)
);

FILL FILL410400x59280 (
);

FILL FILL236360x291460 (
);

OR2X2 _9673_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .B(_662__bF$buf0),
    .Y(_634_)
);

OR2X2 _9253_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .B(_464__bF$buf2),
    .Y(_414_)
);

FILL FILL_0__10914_ (
);

FILL FILL_1__14393_ (
);

NOR2X1 _18956_ (
    .A(_6310__bF$buf2),
    .B(_7857_),
    .Y(_7858_)
);

OR2X2 _18536_ (
    .A(_7440_),
    .B(_7443_),
    .Y(_7444_)
);

OR2X2 _18116_ (
    .A(_7029_),
    .B(_7030_),
    .Y(_7031_)
);

FILL FILL_0__13386_ (
);

AND2X2 _13671_ (
    .A(_3087__bF$buf0),
    .B(\datapath_1.ALUResult [11]),
    .Y(_3155_)
);

MUX2X1 _13251_ (
    .A(_2593_),
    .B(_2548_),
    .S(_2436_),
    .Y(_2796_)
);

FILL FILL_1_BUFX2_insert1105 (
);

FILL FILL_1_BUFX2_insert1107 (
);

FILL FILL_1_BUFX2_insert1109 (
);

FILL FILL286520x306280 (
);

FILL FILL428640x340860 (
);

FILL FILL272840x330980 (
);

FILL FILL_0__9713_ (
);

FILL FILL107920x242060 (
);

FILL FILL412680x54340 (
);

DFFSR _14876_ (
    .CLK(clk_bF$buf77),
    .D(_3870_[24]),
    .Q(_2_[24]),
    .R(rst_bF$buf63),
    .S(vdd)
);

OR2X2 _14456_ (
    .A(vdd),
    .B(\datapath_1.Data [29]),
    .Y(_3730_)
);

OR2X2 _14036_ (
    .A(_3450_),
    .B(_3447_),
    .Y(\datapath_1.alu_1.ALUInB [16])
);

FILL FILL285000x64220 (
);

FILL FILL_0__15952_ (
);

FILL FILL_0__15532_ (
);

FILL FILL_0__15112_ (
);

FILL FILL321480x29640 (
);

FILL FILL_1__11098_ (
);

FILL FILL176320x345800 (
);

AND2X2 _10796_ (
    .A(_1202_),
    .B(_1201_),
    .Y(_1191_[5])
);

DFFSR _10376_ (
    .CLK(clk_bF$buf97),
    .D(_927_[17]),
    .Q(\datapath_1.regfile_1.regOut[15] [17]),
    .R(rst_bF$buf84),
    .S(vdd)
);

FILL FILL110960x182780 (
);

FILL FILL_0__16737_ (
);

AND2X2 _16602_ (
    .A(_4217__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_5539_)
);

FILL FILL_0__11872_ (
);

OR2X2 _19494_ (
    .A(gnd),
    .B(_8385__bF$buf2),
    .Y(_8365_)
);

AND2X2 _19074_ (
    .A(_6238__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_7974_)
);

FILL FILL15960x64220 (
);

FILL FILL32680x14820 (
);

FILL FILL316920x207480 (
);

DFFSR _8944_ (
    .CLK(clk_bF$buf82),
    .D(_201_[4]),
    .Q(\datapath_1.regfile_1.regOut[4] [4]),
    .R(rst_bF$buf94),
    .S(vdd)
);

OR2X2 _8524_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .B(_68__bF$buf0),
    .Y(_48_)
);

FILL FILL_1__18529_ (
);

FILL FILL_1__13244_ (
);

FILL FILL124640x83980 (
);

OR2X2 _17807_ (
    .A(_6724_),
    .B(_6725_),
    .Y(_6726_)
);

FILL FILL16720x217360 (
);

OAI21X1 _12942_ (
    .A(_2165_),
    .B(_2376__bF$buf3),
    .C(_2505_),
    .Y(_2506_)
);

FILL FILL_0__12237_ (
);

NOR3X1 _12522_ (
    .A(_2110_),
    .B(\control_1.op [3]),
    .C(_2111_),
    .Y(_2112_)
);

OR2X2 _12102_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_1873_)
);

FILL FILL_1_BUFX2_insert725 (
);

FILL FILL_1_BUFX2_insert727 (
);

FILL FILL_1_BUFX2_insert729 (
);

FILL FILL101080x83980 (
);

DFFSR _9729_ (
    .CLK(clk_bF$buf90),
    .D(_597_[15]),
    .Q(\datapath_1.regfile_1.regOut[10] [15]),
    .R(rst_bF$buf108),
    .S(vdd)
);

OR2X2 _9309_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_451_)
);

FILL FILL_0__16490_ (
);

AND2X2 _13727_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [19]),
    .Y(_3203_)
);

FILL FILL221920x14820 (
);

XOR2X1 _13307_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2848_)
);

FILL FILL196080x133380 (
);

FILL FILL472720x59280 (
);

FILL FILL_1__15810_ (
);

FILL FILL251560x350740 (
);

OR2X2 _16199_ (
    .A(_5141_),
    .B(_5140_),
    .Y(_5142_)
);

FILL FILL_0__14803_ (
);

FILL FILL232560x187720 (
);

AND2X2 _17980_ (
    .A(_6229__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_6897_)
);

OR2X2 _17560_ (
    .A(_6479_),
    .B(_6482_),
    .Y(_6483_)
);

FILL FILL_0__17275_ (
);

AND2X2 _17140_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_6069_)
);

FILL FILL_1__10789_ (
);

DFFSR _9482_ (
    .CLK(clk_bF$buf86),
    .D(_465_[26]),
    .Q(\datapath_1.regfile_1.regOut[8] [26]),
    .R(rst_bF$buf27),
    .S(vdd)
);

AND2X2 _9062_ (
    .A(_326_),
    .B(_325_),
    .Y(_267_[29])
);

FILL FILL255360x271700 (
);

FILL FILL_1__19487_ (
);

FILL FILL69920x123500 (
);

FILL FILL_0__10303_ (
);

AND2X2 _18765_ (
    .A(_6297__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_7670_)
);

AND2X2 _18345_ (
    .A(_6264__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_7256_)
);

FILL FILL_0__13195_ (
);

OR2X2 _13480_ (
    .A(\datapath_1.PCJump [15]),
    .B(_3005_),
    .Y(_3010_)
);

AND2X2 _13060_ (
    .A(_2616_),
    .B(_2469_),
    .Y(_2617_)
);

FILL FILL_0__19421_ (
);

FILL FILL_0__19001_ (
);

FILL FILL386840x350740 (
);

FILL FILL492480x103740 (
);

FILL FILL_1__12515_ (
);

FILL FILL304000x350740 (
);

FILL FILL_0__9942_ (
);

FILL FILL_0__11508_ (
);

FILL FILL_0__9102_ (
);

FILL FILL313120x54340 (
);

FILL FILL505400x103740 (
);

FILL FILL86640x360620 (
);

OR2X2 _14685_ (
    .A(\datapath_1.rd1 [19]),
    .B(_3869__bF$buf4),
    .Y(_3843_)
);

OR2X2 _14265_ (
    .A(\datapath_1.ALUResult [8]),
    .B(_3671__bF$buf4),
    .Y(_3623_)
);

FILL FILL67640x197600 (
);

FILL FILL294120x4940 (
);

FILL FILL434720x0 (
);

FILL FILL_0__15761_ (
);

FILL FILL_0__15341_ (
);

FILL FILL152000x261820 (
);

FILL FILL_1__17553_ (
);

OR2X2 _10185_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_895_)
);

FILL FILL_1__17133_ (
);

FILL FILL186960x83980 (
);

AND2X2 _16831_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_5764_)
);

FILL FILL_0__16126_ (
);

AND2X2 _16411_ (
    .A(_4210__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_5351_)
);

FILL FILL370880x83980 (
);

FILL FILL40280x207480 (
);

FILL FILL_0__11681_ (
);

FILL FILL_0__11261_ (
);

FILL FILL230280x370500 (
);

AND2X2 _8753_ (
    .A(_160_),
    .B(_159_),
    .Y(_135_[12])
);

FILL FILL_1__13893_ (
);

INVX1 _17616_ (
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_6538_)
);

FILL FILL297920x301340 (
);

FILL FILL367080x202540 (
);

AND2X2 _12751_ (
    .A(_2303_),
    .B(_2315_),
    .Y(_2316_)
);

FILL FILL_0__12466_ (
);

OR2X2 _12331_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .B(_2048__bF$buf0),
    .Y(_1986_)
);

OR2X2 _9958_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .B(_794__bF$buf0),
    .Y(_784_)
);

OR2X2 _9538_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .B(_596__bF$buf4),
    .Y(_564_)
);

OR2X2 _9118_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .B(_398__bF$buf3),
    .Y(_344_)
);

FILL FILL61560x138320 (
);

FILL FILL164160x296400 (
);

FILL FILL121600x192660 (
);

FILL FILL_0_BUFX2_insert380 (
);

FILL FILL42560x296400 (
);

FILL FILL_0_BUFX2_insert382 (
);

AND2X2 _13956_ (
    .A(_3350__bF$buf0),
    .B(_2_[5]),
    .Y(_3382_)
);

FILL FILL_0_BUFX2_insert384 (
);

AND2X2 _13536_ (
    .A(_3045_),
    .B(_3044_),
    .Y(_1_[15])
);

AND2X2 _13116_ (
    .A(_2668_),
    .B(_2297_),
    .Y(_2669_)
);

FILL FILL_0_BUFX2_insert386 (
);

FILL FILL_0_BUFX2_insert388 (
);

FILL FILL_0_BUFX2_insert389 (
);

FILL FILL10640x9880 (
);

FILL FILL196080x271700 (
);

FILL FILL_0__17084_ (
);

FILL FILL382280x286520 (
);

OR2X2 _9291_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_439_)
);

FILL FILL505400x330980 (
);

FILL FILL22040x182780 (
);

FILL FILL_0__15817_ (
);

FILL FILL_0__10952_ (
);

AND2X2 _18994_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_7895_)
);

OR2X2 _18574_ (
    .A(_7481_),
    .B(_7480_),
    .Y(_7482_)
);

OR2X2 _18154_ (
    .A(_7067_),
    .B(_7054_),
    .Y(_7068_)
);

FILL FILL491720x29640 (
);

FILL FILL281200x202540 (
);

FILL FILL_1__12744_ (
);

FILL FILL308560x266760 (
);

FILL FILL_0__9751_ (
);

FILL FILL_0__11737_ (
);

FILL FILL_0__11317_ (
);

OR2X2 _11602_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .B(_1652__bF$buf4),
    .Y(_1620_)
);

OR2X2 _19359_ (
    .A(_8221_),
    .B(_8254_),
    .Y(_8255_)
);

DFFSR _14494_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[29]),
    .Q(\datapath_1.Data [29]),
    .R(rst_bF$buf85),
    .S(vdd)
);

OR2X2 _14074_ (
    .A(_3481_),
    .B(_3482_),
    .Y(_3483_)
);

OR2X2 _8809_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .B(_200__bF$buf2),
    .Y(_198_)
);

FILL FILL_0__15990_ (
);

FILL FILL175560x340860 (
);

FILL FILL_1__13109_ (
);

XOR2X1 _12807_ (
    .A(_2160_),
    .B(_2371_),
    .Y(_2372_)
);

OR2X2 _15699_ (
    .A(_4649_),
    .B(_4648_),
    .Y(_4650_)
);

AND2X2 _15279_ (
    .A(_4236__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_4237_)
);

FILL FILL_1__17782_ (
);

FILL FILL_0__16775_ (
);

OR2X2 _16640_ (
    .A(_5575_),
    .B(_5574_),
    .Y(_5576_)
);

FILL FILL_0__16355_ (
);

OR2X2 _16220_ (
    .A(_5161_),
    .B(_5162_),
    .Y(_5163_)
);

FILL FILL_0__11490_ (
);

FILL FILL250800x133380 (
);

FILL FILL_0__11070_ (
);

OR2X2 _8982_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_273_)
);

DFFSR _8562_ (
    .CLK(clk_bF$buf89),
    .D(_3_[9]),
    .Q(\datapath_1.regfile_1.regOut[1] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

FILL FILL70680x256880 (
);

FILL FILL205200x256880 (
);

OR2X2 _11199_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_1411_)
);

FILL FILL374680x167960 (
);

OR2X2 _17845_ (
    .A(_6763_),
    .B(_6760_),
    .Y(_6764_)
);

OR2X2 _17425_ (
    .A(_6349_),
    .B(_6342_),
    .Y(_6350_)
);

AND2X2 _17005_ (
    .A(_4197__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_5936_)
);

FILL FILL_0__12695_ (
);

OR2X2 _12980_ (
    .A(_2336_),
    .B(_2317_),
    .Y(_2541_)
);

FILL FILL_0__12275_ (
);

INVX1 _12560_ (
    .A(\control_1.op [3]),
    .Y(_2081_)
);

AND2X2 _12140_ (
    .A(_1898_),
    .B(_1897_),
    .Y(_1851_[23])
);

FILL FILL_0__18921_ (
);

FILL FILL219640x217360 (
);

FILL FILL_0__18501_ (
);

AND2X2 _9767_ (
    .A(_676_),
    .B(_675_),
    .Y(_663_[6])
);

DFFSR _9347_ (
    .CLK(clk_bF$buf95),
    .D(_399_[20]),
    .Q(\datapath_1.regfile_1.regOut[7] [20]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL_1__14067_ (
);

OR2X2 _13765_ (
    .A(_3235_),
    .B(_3232_),
    .Y(\datapath_1.mux_pcsrc.dout [24])
);

NOR2X1 _13345_ (
    .A(_2884_),
    .B(_2881_),
    .Y(_2885_)
);

FILL FILL105640x335920 (
);

FILL FILL_0__14421_ (
);

FILL FILL_0__14001_ (
);

FILL FILL131480x276640 (
);

FILL FILL120840x59280 (
);

FILL FILL_1__16633_ (
);

FILL FILL_0__15626_ (
);

OR2X2 _15911_ (
    .A(_4855_),
    .B(_4858_),
    .Y(_4859_)
);

FILL FILL_0__15206_ (
);

FILL FILL355680x113620 (
);

FILL FILL_0__18098_ (
);

OR2X2 _18383_ (
    .A(_7262_),
    .B(_7293_),
    .Y(_7294_)
);

FILL FILL285760x118560 (
);

FILL FILL_0__9560_ (
);

FILL FILL_0__11966_ (
);

FILL FILL_0__9140_ (
);

AND2X2 _11831_ (
    .A(_1732_),
    .B(_1731_),
    .Y(_1719_[6])
);

DFFSR _11411_ (
    .CLK(clk_bF$buf100),
    .D(_1455_[20]),
    .Q(\datapath_1.regfile_1.regOut[23] [20]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL_0__11126_ (
);

OR2X2 _19168_ (
    .A(_8065_),
    .B(_8064_),
    .Y(_8066_)
);

AND2X2 _8618_ (
    .A(_90_),
    .B(_89_),
    .Y(_69_[10])
);

FILL FILL289560x360620 (
);

FILL FILL_1__13758_ (
);

AND2X2 _12616_ (
    .A(_2180_),
    .B(_2176_),
    .Y(_2181_)
);

FILL FILL34200x207480 (
);

FILL FILL421040x108680 (
);

FILL FILL316160x19760 (
);

AND2X2 _15088_ (
    .A(_4070_),
    .B(_4072_),
    .Y(_4073_)
);

FILL FILL15200x365560 (
);

FILL FILL_0__16584_ (
);

FILL FILL321480x321100 (
);

OR2X2 _8791_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_200__bF$buf4),
    .Y(_186_)
);

FILL FILL371640x98800 (
);

FILL FILL29640x326040 (
);

FILL FILL19000x286520 (
);

FILL FILL260680x217360 (
);

FILL FILL_0__17789_ (
);

OR2X2 _17654_ (
    .A(_6574_),
    .B(_6575_),
    .Y(_6576_)
);

AND2X2 _17234_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_6161_)
);

FILL FILL_0__12084_ (
);

FILL FILL433960x237120 (
);

FILL FILL177840x227240 (
);

FILL FILL423320x197600 (
);

DFFSR _9996_ (
    .CLK(clk_bF$buf96),
    .D(_729_[24]),
    .Q(\datapath_1.regfile_1.regOut[12] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

OR2X2 _9576_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_589_)
);

OR2X2 _9156_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_369_)
);

FILL FILL_0__10817_ (
);

FILL FILL_0_BUFX2_insert760 (
);

OR2X2 _18859_ (
    .A(_7760_),
    .B(_7761_),
    .Y(_7762_)
);

AND2X2 _18439_ (
    .A(_6272__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_7349_)
);

FILL FILL87400x113620 (
);

FILL FILL_0_BUFX2_insert762 (
);

AND2X2 _18019_ (
    .A(_6262__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_6935_)
);

OR2X2 _13994_ (
    .A(_3414_),
    .B(_3411_),
    .Y(\datapath_1.alu_1.ALUInB [10])
);

FILL FILL_0_BUFX2_insert764 (
);

FILL FILL_0__13289_ (
);

OR2X2 _13574_ (
    .A(ALUOut[28]),
    .B(_3079__bF$buf3),
    .Y(_3071_)
);

FILL FILL_0_BUFX2_insert766 (
);

NOR3X1 _13154_ (
    .A(_2498_),
    .B(_2704_),
    .C(_2290_),
    .Y(_2705_)
);

FILL FILL_0_BUFX2_insert768 (
);

FILL FILL_0_BUFX2_insert769 (
);

FILL FILL290320x271700 (
);

FILL FILL_0__19515_ (
);

FILL FILL_0__14650_ (
);

FILL FILL287280x222300 (
);

FILL FILL_0__14230_ (
);

FILL FILL_1__12609_ (
);

AND2X2 _14779_ (
    .A(_3885_),
    .B(_3884_),
    .Y(_3870_[7])
);

DFFSR _14359_ (
    .CLK(clk_bF$buf62),
    .D(_3606_[23]),
    .Q(ALUOut[23]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL310840x39520 (
);

FILL FILL_1__16022_ (
);

FILL FILL_0__15855_ (
);

OR2X2 _15720_ (
    .A(_4663_),
    .B(_4670_),
    .Y(_4671_)
);

OR2X2 _15300_ (
    .A(_4255_),
    .B(_4256_),
    .Y(_4257_)
);

FILL FILL_0__10990_ (
);

AND2X2 _18192_ (
    .A(_6216__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_7105_)
);

FILL FILL99560x148200 (
);

FILL FILL_1__17647_ (
);

OR2X2 _10699_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .B(_1190__bF$buf1),
    .Y(_1158_)
);

OR2X2 _10279_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_992__bF$buf4),
    .Y(_938_)
);

AND2X2 _16925_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_5857_)
);

OR2X2 _16505_ (
    .A(_5412_),
    .B(_5443_),
    .Y(_5444_)
);

FILL FILL_0__11355_ (
);

OR2X2 _11640_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_1645_)
);

OR2X2 _11220_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_1425_)
);

OR2X2 _19397_ (
    .A(_8291_),
    .B(_8290_),
    .Y(_8292_)
);

OR2X2 _8847_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_203_)
);

BUFX2 _8427_ (
    .A(_2_[3]),
    .Y(memoryWriteData[3])
);

NAND2X1 _12845_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2410_)
);

DFFSR _12425_ (
    .CLK(clk_bF$buf17),
    .D(_1983_[2]),
    .Q(\datapath_1.regfile_1.regOut[31] [2]),
    .R(rst_bF$buf49),
    .S(vdd)
);

AND2X2 _12005_ (
    .A(_1828_),
    .B(_1827_),
    .Y(_1785_[21])
);

FILL FILL228760x286520 (
);

FILL FILL_0__13501_ (
);

FILL FILL_1__8589_ (
);

FILL FILL_0__16393_ (
);

FILL FILL_1__9950_ (
);

FILL FILL161880x39520 (
);

FILL FILL_0__14706_ (
);

AND2X2 _17883_ (
    .A(_6229__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_6801_)
);

FILL FILL_0__17598_ (
);

OR2X2 _17463_ (
    .A(_6387_),
    .B(_6384_),
    .Y(_6388_)
);

FILL FILL_0__17178_ (
);

OR2X2 _17043_ (
    .A(_5971_),
    .B(_5972_),
    .Y(_5973_)
);

FILL FILL74480x247000 (
);

FILL FILL397480x321100 (
);

FILL FILL209000x247000 (
);

FILL FILL336680x49400 (
);

OR2X2 _9385_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .B(_530__bF$buf0),
    .Y(_482_)
);

FILL FILL104880x330980 (
);

FILL FILL_0__8640_ (
);

FILL FILL9880x54340 (
);

OR2X2 _10911_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_1259_)
);

FILL FILL_0__10206_ (
);

AND2X2 _18668_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_7574_)
);

AND2X2 _18248_ (
    .A(_6211__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_7161_)
);

AND2X2 _13383_ (
    .A(_2919_),
    .B(_2171_),
    .Y(_2920_)
);

FILL FILL432440x103740 (
);

FILL FILL_1__12838_ (
);

FILL FILL165680x39520 (
);

FILL FILL_0__9425_ (
);

FILL FILL_0__9005_ (
);

OR2X2 _14588_ (
    .A(IRWrite_bF$buf2),
    .B(\control_1.op [4]),
    .Y(_3798_)
);

OR2X2 _14168_ (
    .A(\datapath_1.Data [8]),
    .B(_3605__bF$buf3),
    .Y(_3557_)
);

FILL FILL_1__16251_ (
);

FILL FILL_0__15244_ (
);

FILL FILL430160x177840 (
);

FILL FILL407360x88920 (
);

AND2X2 _10088_ (
    .A(_850_),
    .B(_849_),
    .Y(_795_[27])
);

FILL FILL_0__16869_ (
);

AND2X2 _16734_ (
    .A(_4177__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_5669_)
);

FILL FILL_0__16449_ (
);

FILL FILL_0__16029_ (
);

AND2X2 _16314_ (
    .A(_5255_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd2 [16])
);

FILL FILL60800x286520 (
);

FILL FILL101840x4940 (
);

FILL FILL383800x360620 (
);

FILL FILL200640x281580 (
);

FILL FILL497800x108680 (
);

OR2X2 _8656_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .B(_134__bF$buf4),
    .Y(_116_)
);

AND2X2 _17939_ (
    .A(_6317__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_6856_)
);

OR2X2 _17519_ (
    .A(_6442_),
    .B(_6441_),
    .Y(_6443_)
);

FILL FILL_0__12789_ (
);

FILL FILL_0__12369_ (
);

XNOR2X1 _12654_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2219_)
);

OR2X2 _12234_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_1941_)
);

FILL FILL92720x261820 (
);

FILL FILL199120x34580 (
);

FILL FILL89680x212420 (
);

FILL FILL_0__13730_ (
);

FILL FILL_0__13310_ (
);

FILL FILL237120x207480 (
);

FILL FILL_1__8398_ (
);

FILL FILL_0_BUFX2_insert1111 (
);

FILL FILL_0_BUFX2_insert1112 (
);

FILL FILL_0_BUFX2_insert1113 (
);

FILL FILL_0_BUFX2_insert1114 (
);

FILL FILL_0_BUFX2_insert1115 (
);

FILL FILL_0_BUFX2_insert1117 (
);

FILL FILL_0_BUFX2_insert1119 (
);

FILL FILL18240x281580 (
);

OR2X2 _13859_ (
    .A(\datapath_1.a [14]),
    .B(_3342__bF$buf1),
    .Y(_3306_)
);

AND2X2 _13439_ (
    .A(_2972_),
    .B(_2966_),
    .Y(_2973_)
);

NAND2X1 _13019_ (
    .A(_2329_),
    .B(_2548_),
    .Y(_2578_)
);

FILL FILL_1__15102_ (
);

FILL FILL_0__14935_ (
);

AND2X2 _14800_ (
    .A(_3899_),
    .B(_3898_),
    .Y(_3870_[14])
);

FILL FILL_0__14515_ (
);

FILL FILL280440x158080 (
);

FILL FILL298680x0 (
);

AND2X2 _17692_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_6613_)
);

OR2X2 _17272_ (
    .A(_6198_),
    .B(_6183_),
    .Y(_6199_)
);

FILL FILL421040x49400 (
);

AND2X2 _9194_ (
    .A(_394_),
    .B(_393_),
    .Y(_333_[30])
);

FILL FILL239400x296400 (
);

OR2X2 _10720_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_1190__bF$buf2),
    .Y(_1172_)
);

FILL FILL_0__10435_ (
);

FILL FILL_0__10015_ (
);

OR2X2 _10300_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .B(_992__bF$buf1),
    .Y(_952_)
);

AND2X2 _18897_ (
    .A(_6323__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_7800_)
);

OR2X2 _18477_ (
    .A(_7385_),
    .B(_7384_),
    .Y(_7386_)
);

OR2X2 _18057_ (
    .A(_6972_),
    .B(_6956_),
    .Y(_6973_)
);

AOI21X1 _13192_ (
    .A(_2417_),
    .B(_2740_),
    .C(_2738_),
    .Y(_2741_)
);

FILL FILL_0__19133_ (
);

FILL FILL476520x128440 (
);

DFFSR _11925_ (
    .CLK(clk_bF$buf52),
    .D(_1719_[18]),
    .Q(\datapath_1.regfile_1.regOut[27] [18]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL_0__9234_ (
);

OR2X2 _11505_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_1575_)
);

FILL FILL90440x123500 (
);

OR2X2 _14397_ (
    .A(memoryOutData[9]),
    .B(_3737__bF$buf4),
    .Y(_3691_)
);

FILL FILL_0__15893_ (
);

FILL FILL_0__15473_ (
);

FILL FILL_0__15053_ (
);

FILL FILL115520x340860 (
);

FILL FILL141360x281580 (
);

FILL FILL_0__16678_ (
);

AND2X2 _16963_ (
    .A(_4154__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_5894_)
);

OR2X2 _16543_ (
    .A(_5479_),
    .B(_5480_),
    .Y(_5481_)
);

FILL FILL_0__16258_ (
);

FILL FILL16720x103740 (
);

AND2X2 _16123_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_5067_)
);

FILL FILL132240x256880 (
);

FILL FILL272080x49400 (
);

AND2X2 _8885_ (
    .A(_228_),
    .B(_227_),
    .Y(_201_[13])
);

AND2X2 _8465_ (
    .A(_8_),
    .B(_7_),
    .Y(_3_[2])
);

FILL FILL_1__13185_ (
);

FILL FILL314640x167960 (
);

AND2X2 _17748_ (
    .A(_6236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_6668_)
);

AND2X2 _17328_ (
    .A(_6203_),
    .B(_6227_),
    .Y(_6254_)
);

AND2X2 _12883_ (
    .A(_2440_),
    .B(_2447_),
    .Y(_2448_)
);

FILL FILL_1__19411_ (
);

NAND3X1 _12463_ (
    .A(_2055_),
    .B(_2056_),
    .C(_2053_),
    .Y(_2057_)
);

DFFSR _12043_ (
    .CLK(clk_bF$buf39),
    .D(_1785_[7]),
    .Q(\datapath_1.regfile_1.regOut[28] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

FILL FILL_0__18404_ (
);

FILL FILL_1_BUFX2_insert1070 (
);

FILL FILL363280x192660 (
);

FILL FILL_1_BUFX2_insert1072 (
);

AND2X2 _13668_ (
    .A(_3081__bF$buf1),
    .B(ALUOut[11]),
    .Y(_3152_)
);

FILL FILL37240x261820 (
);

OAI21X1 _13248_ (
    .A(_2790_),
    .B(_2792_),
    .C(_2237_),
    .Y(_2793_)
);

FILL FILL_1__15751_ (
);

FILL FILL455240x148200 (
);

FILL FILL_0__14324_ (
);

OR2X2 _17081_ (
    .A(_6010_),
    .B(_5979_),
    .Y(_6011_)
);

FILL FILL_1__16116_ (
);

FILL FILL_0__15949_ (
);

FILL FILL325280x59280 (
);

AND2X2 _15814_ (
    .A(_4203__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_4763_)
);

FILL FILL_0__15109_ (
);

AND2X2 _18286_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_7198_)
);

FILL FILL_0__19362_ (
);

FILL FILL_1__12876_ (
);

FILL FILL_1__12456_ (
);

FILL FILL417240x207480 (
);

FILL FILL504640x212420 (
);

FILL FILL_0__9883_ (
);

FILL FILL_0__11869_ (
);

FILL FILL_0__11449_ (
);

OR2X2 _11734_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .B(_1718__bF$buf1),
    .Y(_1688_)
);

OR2X2 _11314_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .B(_1520__bF$buf2),
    .Y(_1468_)
);

FILL FILL_0__12810_ (
);

FILL FILL415720x375440 (
);

FILL FILL_1_BUFX2_insert690 (
);

NAND3X1 _12939_ (
    .A(_2386_),
    .B(ALUControl[1]),
    .C(ALUControl[0]),
    .Y(_2503_)
);

FILL FILL_1_BUFX2_insert692 (
);

OAI21X1 _12519_ (
    .A(\control_1.reg_state.dout [2]),
    .B(_2107_),
    .C(_2109_),
    .Y(ALUSrcB[1])
);

FILL FILL_1__17074_ (
);

OR2X2 _16772_ (
    .A(_5704_),
    .B(_5705_),
    .Y(_5706_)
);

FILL FILL_0__16067_ (
);

OR2X2 _16352_ (
    .A(_5292_),
    .B(_5289_),
    .Y(_5293_)
);

DFFSR _8694_ (
    .CLK(clk_bF$buf28),
    .D(_69_[12]),
    .Q(\datapath_1.regfile_1.regOut[2] [12]),
    .R(rst_bF$buf0),
    .S(vdd)
);

FILL FILL269040x360620 (
);

FILL FILL202160x44460 (
);

BUFX2 BUFX2_insert360 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf0 )
);

BUFX2 BUFX2_insert361 (
    .A(_4175_),
    .Y(_4175__bF$buf4)
);

BUFX2 BUFX2_insert362 (
    .A(_4175_),
    .Y(_4175__bF$buf3)
);

BUFX2 BUFX2_insert363 (
    .A(_4175_),
    .Y(_4175__bF$buf2)
);

NOR2X1 _17977_ (
    .A(_6310__bF$buf0),
    .B(_6893_),
    .Y(_6894_)
);

BUFX2 BUFX2_insert364 (
    .A(_4175_),
    .Y(_4175__bF$buf1)
);

AND2X2 _17557_ (
    .A(_6216__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_6480_)
);

BUFX2 BUFX2_insert365 (
    .A(_4175_),
    .Y(_4175__bF$buf0)
);

BUFX2 BUFX2_insert366 (
    .A(_6321_),
    .Y(_6321__bF$buf4)
);

AND2X2 _17137_ (
    .A(_4177__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_6066_)
);

BUFX2 BUFX2_insert367 (
    .A(_6321_),
    .Y(_6321__bF$buf3)
);

BUFX2 BUFX2_insert368 (
    .A(_6321_),
    .Y(_6321__bF$buf2)
);

AND2X2 _12692_ (
    .A(_2251_),
    .B(_2256_),
    .Y(_2257_)
);

BUFX2 BUFX2_insert369 (
    .A(_6321_),
    .Y(_6321__bF$buf1)
);

AND2X2 _12272_ (
    .A(_1966_),
    .B(_1965_),
    .Y(_1917_[24])
);

FILL FILL_0__18633_ (
);

FILL FILL77520x365560 (
);

FILL FILL_0__18213_ (
);

AND2X2 _9899_ (
    .A(_744_),
    .B(_743_),
    .Y(_729_[7])
);

DFFSR _9479_ (
    .CLK(clk_bF$buf73),
    .D(_465_[23]),
    .Q(\datapath_1.regfile_1.regOut[8] [23]),
    .R(rst_bF$buf39),
    .S(vdd)
);

AND2X2 _9059_ (
    .A(_324_),
    .B(_323_),
    .Y(_267_[28])
);

FILL FILL_1__11727_ (
);

FILL FILL_1__14199_ (
);

OR2X2 _13897_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [27]),
    .Y(_3331_)
);

OR2X2 _13477_ (
    .A(\datapath_1.PCJump [14]),
    .B(_3005_),
    .Y(_3008_)
);

OR2X2 _13057_ (
    .A(_2454_),
    .B(_2449_),
    .Y(_2614_)
);

FILL FILL_1__15140_ (
);

FILL FILL229520x44460 (
);

FILL FILL_0__19418_ (
);

FILL FILL_0__14553_ (
);

FILL FILL_0__14133_ (
);

FILL FILL278920x0 (
);

FILL FILL_0__9519_ (
);

FILL FILL323760x79040 (
);

FILL FILL_1__16765_ (
);

FILL FILL_0__15758_ (
);

FILL FILL_0__15338_ (
);

OR2X2 _15623_ (
    .A(_4574_),
    .B(_4573_),
    .Y(_4575_)
);

AND2X2 _15203_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_4161_)
);

FILL FILL_0__10053_ (
);

AND2X2 _18095_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_7010_)
);

FILL FILL288800x306280 (
);

FILL FILL71440x306280 (
);

FILL FILL375440x217360 (
);

AND2X2 _16828_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_5761_)
);

OR2X2 _16408_ (
    .A(_5347_),
    .B(_5340_),
    .Y(_5348_)
);

FILL FILL_0__9692_ (
);

FILL FILL_0__9272_ (
);

AND2X2 _11963_ (
    .A(_1800_),
    .B(_1799_),
    .Y(_1785_[7])
);

FILL FILL_1__18911_ (
);

DFFSR _11543_ (
    .CLK(clk_bF$buf26),
    .D(_1521_[23]),
    .Q(\datapath_1.regfile_1.regOut[24] [23]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL_0__11258_ (
);

AND2X2 _11123_ (
    .A(_1380_),
    .B(_1379_),
    .Y(_1323_[28])
);

FILL FILL_0__15091_ (
);

FILL FILL379240x138320 (
);

NAND2X1 _12748_ (
    .A(\datapath_1.alu_1.ALUInA [23]),
    .B(_2312_),
    .Y(_2313_)
);

FILL FILL178600x345800 (
);

OR2X2 _12328_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(_2048__bF$buf0),
    .Y(_1984_)
);

FILL FILL_1__14831_ (
);

FILL FILL_0__13824_ (
);

FILL FILL101080x340860 (
);

AND2X2 _16581_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_5518_)
);

FILL FILL_0__16296_ (
);

AND2X2 _16161_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_5105_)
);

FILL FILL38760x64220 (
);

FILL FILL415720x24700 (
);

FILL FILL291080x197600 (
);

FILL FILL_1__15616_ (
);

FILL FILL_1__18088_ (
);

FILL FILL459040x69160 (
);

AND2X2 _17786_ (
    .A(_6216__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_6706_)
);

OR2X2 _17366_ (
    .A(_6286_),
    .B(_6291_),
    .Y(_6292_)
);

OR2X2 _12081_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_1859_)
);

FILL FILL367840x232180 (
);

FILL FILL_0__18862_ (
);

FILL FILL_0__18442_ (
);

FILL FILL_0__18022_ (
);

OR2X2 _9288_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_437_)
);

FILL FILL267520x326040 (
);

FILL FILL_0__8543_ (
);

FILL FILL_0__10949_ (
);

AND2X2 _10814_ (
    .A(_1214_),
    .B(_1213_),
    .Y(_1191_[11])
);

FILL FILL_0__10529_ (
);

FILL FILL253840x350740 (
);

NOR2X1 _13286_ (
    .A(_2210_),
    .B(_2425_),
    .Y(_2829_)
);

OR2X2 _19512_ (
    .A(gnd),
    .B(_8385__bF$buf2),
    .Y(_8377_)
);

FILL FILL_0__19227_ (
);

FILL FILL419520x24700 (
);

FILL FILL_0__14782_ (
);

FILL FILL253080x256880 (
);

FILL FILL79040x29640 (
);

FILL FILL257640x271700 (
);

FILL FILL11400x143260 (
);

FILL FILL15200x49400 (
);

FILL FILL_1__16574_ (
);

AND2X2 _15852_ (
    .A(_4228__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_4801_)
);

FILL FILL_0__15567_ (
);

FILL FILL_0__15147_ (
);

OR2X2 _15432_ (
    .A(_4383_),
    .B(_4386_),
    .Y(_4387_)
);

DFFSR _15012_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[31]),
    .Q(\datapath_1.PCJump [31]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL161120x44460 (
);

FILL FILL494760x103740 (
);

FILL FILL351120x133380 (
);

OR2X2 _16637_ (
    .A(_5571_),
    .B(_5572_),
    .Y(_5573_)
);

FILL FILL403560x301340 (
);

OR2X2 _16217_ (
    .A(_5159_),
    .B(_5144_),
    .Y(_5160_)
);

FILL FILL211280x118560 (
);

OR2X2 _11772_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_1713_)
);

OR2X2 _11352_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_1493_)
);

FILL FILL_0__11067_ (
);

FILL FILL_0__17713_ (
);

OR2X2 _8979_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_271_)
);

DFFSR _8559_ (
    .CLK(clk_bF$buf59),
    .D(_3_[6]),
    .Q(\datapath_1.regfile_1.regOut[1] [6]),
    .R(rst_bF$buf106),
    .S(vdd)
);

FILL FILL173280x232180 (
);

FILL FILL148960x0 (
);

FILL FILL410400x271700 (
);

AND2X2 _9920_ (
    .A(_758_),
    .B(_757_),
    .Y(_729_[14])
);

AND2X2 _9500_ (
    .A(_538_),
    .B(_537_),
    .Y(_531_[3])
);

FILL FILL_1__13699_ (
);

FILL FILL372400x44460 (
);

FILL FILL_1__13279_ (
);

FILL FILL145920x138320 (
);

INVX1 _12977_ (
    .A(_2538_),
    .Y(\datapath_1.ALUResult [28])
);

AND2X2 _12557_ (
    .A(_2110_),
    .B(\control_1.op [3]),
    .Y(_2078_)
);

AND2X2 _12137_ (
    .A(_1896_),
    .B(_1895_),
    .Y(_1851_[22])
);

FILL FILL_1__14640_ (
);

FILL FILL_0__18918_ (
);

FILL FILL505400x177840 (
);

FILL FILL_0__13213_ (
);

FILL FILL19000x172900 (
);

FILL FILL145160x365560 (
);

FILL FILL232560x370500 (
);

AND2X2 _16390_ (
    .A(_4187__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_5330_)
);

FILL FILL346560x118560 (
);

FILL FILL4560x301340 (
);

FILL FILL_1__10980_ (
);

FILL FILL_0__14838_ (
);

FILL FILL369360x202540 (
);

OR2X2 _14703_ (
    .A(\datapath_1.rd1 [25]),
    .B(_3869__bF$buf4),
    .Y(_3855_)
);

BUFX2 BUFX2_insert740 (
    .A(_4239_),
    .Y(_4239__bF$buf3)
);

BUFX2 BUFX2_insert741 (
    .A(_4239_),
    .Y(_4239__bF$buf2)
);

BUFX2 BUFX2_insert742 (
    .A(_4239_),
    .Y(_4239__bF$buf1)
);

BUFX2 BUFX2_insert743 (
    .A(_4239_),
    .Y(_4239__bF$buf0)
);

FILL FILL82840x301340 (
);

BUFX2 BUFX2_insert744 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf3 )
);

FILL FILL106400x182780 (
);

AND2X2 _17595_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_6518_)
);

BUFX2 BUFX2_insert745 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf2 )
);

BUFX2 BUFX2_insert746 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf1 )
);

OR2X2 _17175_ (
    .A(_6099_),
    .B(_6102_),
    .Y(_6103_)
);

BUFX2 BUFX2_insert747 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf0 )
);

BUFX2 BUFX2_insert748 (
    .A(_1520_),
    .Y(_1520__bF$buf4)
);

BUFX2 BUFX2_insert749 (
    .A(_1520_),
    .Y(_1520__bF$buf3)
);

FILL FILL63840x138320 (
);

FILL FILL69160x212420 (
);

FILL FILL_0__18671_ (
);

FILL FILL490200x148200 (
);

FILL FILL431680x98800 (
);

FILL FILL243200x242060 (
);

FILL FILL82080x207480 (
);

DFFSR _9097_ (
    .CLK(clk_bF$buf67),
    .D(_267_[28]),
    .Q(\datapath_1.regfile_1.regOut[5] [28]),
    .R(rst_bF$buf7),
    .S(vdd)
);

FILL FILL_1__11345_ (
);

AND2X2 _15908_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_4856_)
);

FILL FILL437760x4940 (
);

FILL FILL_0__8772_ (
);

FILL FILL_0__10338_ (
);

DFFSR _10623_ (
    .CLK(clk_bF$buf29),
    .D(_1059_[6]),
    .Q(\datapath_1.regfile_1.regOut[17] [6]),
    .R(rst_bF$buf48),
    .S(vdd)
);

OR2X2 _10203_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_907_)
);

NAND3X1 _13095_ (
    .A(_2602_),
    .B(_2307_),
    .C(_2524_),
    .Y(_2650_)
);

FILL FILL77520x49400 (
);

FILL FILL_0__19456_ (
);

FILL FILL247000x163020 (
);

AND2X2 _19321_ (
    .A(_6264__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_8217_)
);

FILL FILL_0__14171_ (
);

FILL FILL384560x286520 (
);

FILL FILL_0__9137_ (
);

AND2X2 _11828_ (
    .A(_1730_),
    .B(_1729_),
    .Y(_1719_[5])
);

DFFSR _11408_ (
    .CLK(clk_bF$buf76),
    .D(_1455_[17]),
    .Q(\datapath_1.regfile_1.regOut[23] [17]),
    .R(rst_bF$buf112),
    .S(vdd)
);

FILL FILL_0__15796_ (
);

FILL FILL_0__15376_ (
);

AND2X2 _15661_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_4613_)
);

OR2X2 _15241_ (
    .A(_4198_),
    .B(_4196_),
    .Y(_4199_)
);

FILL FILL41800x192660 (
);

FILL FILL_0__10091_ (
);

FILL FILL_1__8933_ (
);

FILL FILL334400x74100 (
);

FILL FILL433200x365560 (
);

FILL FILL_1__17588_ (
);

AND2X2 _16866_ (
    .A(_4210__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_5799_)
);

AND2X2 _16446_ (
    .A(_4181__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_5385_)
);

AND2X2 _16026_ (
    .A(_4175__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_4972_)
);

OR2X2 _11581_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .B(_1652__bF$buf0),
    .Y(_1606_)
);

FILL FILL_0__11296_ (
);

DFFSR _11161_ (
    .CLK(clk_bF$buf52),
    .D(_1323_[28]),
    .Q(\datapath_1.regfile_1.regOut[21] [28]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL278920x321100 (
);

FILL FILL25080x148200 (
);

FILL FILL348080x222300 (
);

FILL FILL_0__17522_ (
);

FILL FILL437000x286520 (
);

FILL FILL_0__17102_ (
);

OR2X2 _8788_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .B(_200__bF$buf0),
    .Y(_184_)
);

FILL FILL_1__10616_ (
);

FILL FILL180120x14820 (
);

INVX1 _12786_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .Y(_2351_)
);

OR2X2 _12366_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_2009_)
);

FILL FILL_0__18727_ (
);

FILL FILL_0__18307_ (
);

FILL FILL112480x158080 (
);

FILL FILL_0__13862_ (
);

FILL FILL_0__13442_ (
);

FILL FILL_0__8408_ (
);

FILL FILL_1__9891_ (
);

FILL FILL72960x256880 (
);

FILL FILL78280x330980 (
);

FILL FILL_1__15234_ (
);

AND2X2 _14932_ (
    .A(_3967_),
    .B(_3966_),
    .Y(_3936_[15])
);

AND2X2 _14512_ (
    .A(_3747_),
    .B(_3746_),
    .Y(_3738_[4])
);

FILL FILL330600x340860 (
);

FILL FILL_0__18480_ (
);

FILL FILL_0__18060_ (
);

FILL FILL_1__16439_ (
);

AND2X2 _15717_ (
    .A(_4210__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_4668_)
);

FILL FILL139840x123500 (
);

FILL FILL107160x69160 (
);

FILL FILL_0__10987_ (
);

FILL FILL_0__10567_ (
);

OR2X2 _10852_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .B(_1256__bF$buf2),
    .Y(_1240_)
);

OR2X2 _10432_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .B(_1058__bF$buf3),
    .Y(_1020_)
);

FILL FILL_0__10147_ (
);

OR2X2 _10012_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .B(_860__bF$buf3),
    .Y(_800_)
);

OR2X2 _18189_ (
    .A(_7068_),
    .B(_7102_),
    .Y(_7103_)
);

DFFSR _19550_ (
    .CLK(clk_bF$buf14),
    .D(_8320_[27]),
    .Q(\datapath_1.regfile_1.regOut[0] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

AND2X2 _19130_ (
    .A(_6282__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_8029_)
);

FILL FILL429400x167960 (
);

OR2X2 _11637_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_1643_)
);

OR2X2 _11217_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_1423_)
);

FILL FILL_1__13720_ (
);

FILL FILL357960x113620 (
);

FILL FILL_0__12713_ (
);

FILL FILL_1__16192_ (
);

AND2X2 _15890_ (
    .A(_4225__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_4838_)
);

OR2X2 _15470_ (
    .A(_4424_),
    .B(_4423_),
    .Y(_4425_)
);

FILL FILL_0__15185_ (
);

OAI21X1 _15050_ (
    .A(_4038_),
    .B(_4007_),
    .C(_4017_),
    .Y(_4039_)
);

FILL FILL_1__14925_ (
);

FILL FILL_0__13918_ (
);

FILL FILL167200x232180 (
);

OR2X2 _16675_ (
    .A(_5610_),
    .B(_5609_),
    .Y(_5611_)
);

AND2X2 _16255_ (
    .A(_4225__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_5197_)
);

AND2X2 _11390_ (
    .A(_1518_),
    .B(_1517_),
    .Y(_1455_[31])
);

FILL FILL_1__9107_ (
);

FILL FILL_0__17751_ (
);

FILL FILL_0__17331_ (
);

AND2X2 _8597_ (
    .A(_76_),
    .B(_75_),
    .Y(_69_[3])
);

FILL FILL_1__10425_ (
);

FILL FILL55480x197600 (
);

FILL FILL423320x108680 (
);

FILL FILL254600x103740 (
);

NAND2X1 _12595_ (
    .A(_2158_),
    .B(_2159_),
    .Y(_2160_)
);

DFFSR _12175_ (
    .CLK(clk_bF$buf107),
    .D(_1851_[10]),
    .Q(\datapath_1.regfile_1.regOut[29] [10]),
    .R(rst_bF$buf88),
    .S(vdd)
);

FILL FILL49400x153140 (
);

FILL FILL_0__18956_ (
);

OR2X2 _18821_ (
    .A(_7717_),
    .B(_7724_),
    .Y(_7725_)
);

FILL FILL_0__18536_ (
);

AND2X2 _18401_ (
    .A(_6315__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_7311_)
);

FILL FILL_0__13671_ (
);

FILL FILL_0__13251_ (
);

FILL FILL466640x34580 (
);

INVX2 _10908_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .Y(_1322_)
);

FILL FILL262960x217360 (
);

DFFSR _14741_ (
    .CLK(clk_bF$buf38),
    .D(_3804_[18]),
    .Q(\datapath_1.a [18]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL_0__14456_ (
);

FILL FILL_0__14036_ (
);

OR2X2 _14321_ (
    .A(vdd),
    .B(ALUOut[27]),
    .Y(_3660_)
);

FILL FILL504640x49400 (
);

FILL FILL_1__16668_ (
);

AND2X2 _15946_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_4893_)
);

OR2X2 _15526_ (
    .A(_4479_),
    .B(_4478_),
    .Y(_4480_)
);

AND2X2 _15106_ (
    .A(_4039_),
    .B(_4084_),
    .Y(_4087_)
);

FILL FILL_0__8390_ (
);

FILL FILL_0__10796_ (
);

AND2X2 _10661_ (
    .A(_1132_),
    .B(_1131_),
    .Y(_1125_[3])
);

DFFSR _10241_ (
    .CLK(clk_bF$buf71),
    .D(_861_[11]),
    .Q(\datapath_1.regfile_1.regOut[14] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL292600x271700 (
);

FILL FILL_0__16602_ (
);

FILL FILL_0__19494_ (
);

FILL FILL_0__19074_ (
);

OR2X2 _11866_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_1784__bF$buf3),
    .Y(_1756_)
);

FILL FILL_0__9175_ (
);

FILL FILL344280x345800 (
);

OR2X2 _11446_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_1586__bF$buf1),
    .Y(_1536_)
);

DFFSR _11026_ (
    .CLK(clk_bF$buf84),
    .D(_1257_[22]),
    .Q(\datapath_1.regfile_1.regOut[20] [22]),
    .R(rst_bF$buf47),
    .S(vdd)
);

FILL FILL_0__17807_ (
);

FILL FILL_0__12942_ (
);

FILL FILL_0__12522_ (
);

FILL FILL233320x123500 (
);

FILL FILL_0__13727_ (
);

FILL FILL_0__13307_ (
);

FILL FILL_0_BUFX2_insert1080 (
);

FILL FILL_0_BUFX2_insert1082 (
);

AND2X2 _16484_ (
    .A(_4167__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_5423_)
);

FILL FILL_0__16199_ (
);

OR2X2 _16064_ (
    .A(_5008_),
    .B(_5007_),
    .Y(_5009_)
);

FILL FILL_0_BUFX2_insert1084 (
);

FILL FILL_0_BUFX2_insert1086 (
);

FILL FILL_0_BUFX2_insert1087 (
);

FILL FILL_0_BUFX2_insert1088 (
);

FILL FILL_0_BUFX2_insert1089 (
);

FILL FILL_0__17980_ (
);

FILL FILL_0__17560_ (
);

FILL FILL_0__17140_ (
);

FILL FILL264480x321100 (
);

AND2X2 _17689_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_6610_)
);

OR2X2 _17269_ (
    .A(_6194_),
    .B(_6195_),
    .Y(_6196_)
);

FILL FILL_1__19352_ (
);

FILL FILL194560x326040 (
);

AND2X2 _18630_ (
    .A(_6250__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_7537_)
);

OR2X2 _18210_ (
    .A(_7119_),
    .B(_7122_),
    .Y(_7123_)
);

FILL FILL_0__13060_ (
);

FILL FILL_1__11439_ (
);

FILL FILL_0__8866_ (
);

OR2X2 _10717_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_1190__bF$buf0),
    .Y(_1170_)
);

FILL FILL461320x69160 (
);

OAI21X1 _13189_ (
    .A(_2417_),
    .B(_2376__bF$buf0),
    .C(_2737_),
    .Y(_2738_)
);

FILL FILL_1__15692_ (
);

FILL FILL275880x256880 (
);

AND2X2 _19415_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_8310_)
);

FILL FILL_0__14685_ (
);

OR2X2 _14970_ (
    .A(\datapath_1.mux_pcsrc.dout [28]),
    .B(_4001__bF$buf4),
    .Y(_3993_)
);

FILL FILL_0__14265_ (
);

OR2X2 _14550_ (
    .A(memoryOutData[17]),
    .B(_3803__bF$buf2),
    .Y(_3773_)
);

OR2X2 _14130_ (
    .A(_3529_),
    .B(_3530_),
    .Y(_3531_)
);

FILL FILL376200x335920 (
);

FILL FILL399760x321100 (
);

FILL FILL_1__16057_ (
);

FILL FILL25840x98800 (
);

AND2X2 _15755_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_4705_)
);

OR2X2 _15335_ (
    .A(_4288_),
    .B(_4291_),
    .Y(_4292_)
);

DFFSR _10890_ (
    .CLK(clk_bF$buf90),
    .D(_1191_[15]),
    .Q(\datapath_1.regfile_1.regOut[19] [15]),
    .R(rst_bF$buf108),
    .S(vdd)
);

OR2X2 _10470_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_1045_)
);

FILL FILL_0__10185_ (
);

OR2X2 _10050_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_825_)
);

FILL FILL_0__16831_ (
);

FILL FILL434720x103740 (
);

DFFSR _11675_ (
    .CLK(clk_bF$buf86),
    .D(_1587_[26]),
    .Q(\datapath_1.regfile_1.regOut[25] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

FILL FILL_1__18203_ (
);

AND2X2 _11255_ (
    .A(_1448_),
    .B(_1447_),
    .Y(_1389_[29])
);

AND2X2 _17901_ (
    .A(_6216__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_6819_)
);

FILL FILL_0__12331_ (
);

FILL FILL502360x172900 (
);

OR2X2 _9823_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_728__bF$buf3),
    .Y(_714_)
);

OR2X2 _9403_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_530__bF$buf0),
    .Y(_494_)
);

FILL FILL_1__8780_ (
);

FILL FILL_1__14543_ (
);

FILL FILL_0__13956_ (
);

AND2X2 _13821_ (
    .A(_3280_),
    .B(_3279_),
    .Y(\datapath_1.alu_1.ALUInA [1])
);

FILL FILL_0__13536_ (
);

FILL FILL_0__13116_ (
);

OR2X2 _13401_ (
    .A(_2157__bF$buf1),
    .B(_2936_),
    .Y(_2937_)
);

FILL FILL487160x79040 (
);

AND2X2 _16293_ (
    .A(_4177__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_5235_)
);

DFFSR _14606_ (
    .CLK(clk_bF$buf12),
    .D(_3738_[12]),
    .Q(\datapath_1.PCJump [14]),
    .R(rst_bF$buf91),
    .S(vdd)
);

AND2X2 _17498_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_6422_)
);

OR2X2 _17078_ (
    .A(_6004_),
    .B(_6007_),
    .Y(_6008_)
);

FILL FILL_0__18574_ (
);

FILL FILL294880x370500 (
);

FILL FILL_0__18154_ (
);

FILL FILL_0__8675_ (
);

AND2X2 _10946_ (
    .A(_1282_),
    .B(_1281_),
    .Y(_1257_[12])
);

AND2X2 _10526_ (
    .A(_1062_),
    .B(_1061_),
    .Y(_1059_[1])
);

DFFSR _10106_ (
    .CLK(clk_bF$buf14),
    .D(_795_[5]),
    .Q(\datapath_1.regfile_1.regOut[13] [5]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL_0__11602_ (
);

FILL FILL307040x276640 (
);

FILL FILL282720x158080 (
);

FILL FILL424840x192660 (
);

FILL FILL52440x163020 (
);

FILL FILL_0__19359_ (
);

OR2X2 _19224_ (
    .A(_8120_),
    .B(_8121_),
    .Y(_8122_)
);

FILL FILL_0__12807_ (
);

AND2X2 _15984_ (
    .A(_4225__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_4931_)
);

FILL FILL_0__15279_ (
);

OR2X2 _15564_ (
    .A(_4515_),
    .B(_4516_),
    .Y(_4517_)
);

FILL FILL364040x64220 (
);

NAND2X1 _15144_ (
    .A(_4043_),
    .B(_4080_),
    .Y(_4111_)
);

FILL FILL_0__16640_ (
);

FILL FILL_0__16220_ (
);

FILL FILL277400x375440 (
);

OR2X2 _16769_ (
    .A(_5699_),
    .B(_5702_),
    .Y(_5703_)
);

AND2X2 _16349_ (
    .A(_4158__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_5290_)
);

FILL FILL_1__18852_ (
);

OR2X2 _11484_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_1561_)
);

FILL FILL_0__11199_ (
);

OR2X2 _11064_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_1341_)
);

FILL FILL200640x330980 (
);

FILL FILL_0__17845_ (
);

FILL FILL_0__17425_ (
);

AND2X2 _17710_ (
    .A(_6326__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_6631_)
);

FILL FILL_0__17005_ (
);

FILL FILL_0__12980_ (
);

FILL FILL_0__12560_ (
);

FILL FILL_0__12140_ (
);

AND2X2 _9632_ (
    .A(_606_),
    .B(_605_),
    .Y(_597_[4])
);

DFFSR _9212_ (
    .CLK(clk_bF$buf13),
    .D(_333_[14]),
    .Q(\datapath_1.regfile_1.regOut[6] [14]),
    .R(rst_bF$buf90),
    .S(vdd)
);

INVX1 _12689_ (
    .A(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2254_)
);

FILL FILL_1__19217_ (
);

AND2X2 _12269_ (
    .A(_1964_),
    .B(_1963_),
    .Y(_1917_[23])
);

OR2X2 _18915_ (
    .A(_7815_),
    .B(_7816_),
    .Y(_7817_)
);

FILL FILL_0__13765_ (
);

AND2X2 _13630_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3120_)
);

NAND3X1 _13210_ (
    .A(_2379__bF$buf1),
    .B(\datapath_1.alu_1.ALUInB [14]),
    .C(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2758_)
);

FILL FILL_1__9794_ (
);

FILL FILL322240x148200 (
);

FILL FILL12920x256880 (
);

FILL FILL18240x330980 (
);

FILL FILL_1__15557_ (
);

OR2X2 _14835_ (
    .A(\datapath_1.rd2 [26]),
    .B(_3935__bF$buf2),
    .Y(_3923_)
);

OR2X2 _14415_ (
    .A(memoryOutData[15]),
    .B(_3737__bF$buf4),
    .Y(_3703_)
);

FILL FILL414960x83980 (
);

FILL FILL207480x83980 (
);

FILL FILL_1__11477_ (
);

FILL FILL365560x192660 (
);

DFFSR _10755_ (
    .CLK(clk_bF$buf75),
    .D(_1125_[9]),
    .Q(\datapath_1.regfile_1.regOut[18] [9]),
    .R(rst_bF$buf27),
    .S(vdd)
);

OR2X2 _10335_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_975_)
);

FILL FILL22040x345800 (
);

FILL FILL_0__11831_ (
);

AND2X2 _19453_ (
    .A(_8337_),
    .B(_8336_),
    .Y(_8320_[8])
);

FILL FILL_0__19168_ (
);

OR2X2 _19033_ (
    .A(_7901_),
    .B(_7933_),
    .Y(_7934_)
);

FILL FILL392920x340860 (
);

AND2X2 _8903_ (
    .A(_240_),
    .B(_239_),
    .Y(_201_[19])
);

FILL FILL304760x14820 (
);

FILL FILL_0__9269_ (
);

FILL FILL348080x59280 (
);

FILL FILL_1_BUFX2_insert311 (
);

NOR2X1 _12901_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2466_)
);

FILL FILL_1_BUFX2_insert313 (
);

AND2X2 _15793_ (
    .A(_4175__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_4743_)
);

AND2X2 _15373_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_4329_)
);

FILL FILL386840x0 (
);

OR2X2 _16998_ (
    .A(_5927_),
    .B(_5928_),
    .Y(_5929_)
);

AND2X2 _16578_ (
    .A(_4181__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [21]),
    .Y(_5515_)
);

AND2X2 _16158_ (
    .A(_4146__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_5102_)
);

DFFSR _11293_ (
    .CLK(clk_bF$buf95),
    .D(_1389_[31]),
    .Q(\datapath_1.regfile_1.regOut[22] [31]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL430160x0 (
);

FILL FILL500840x365560 (
);

FILL FILL_0__17654_ (
);

DFFSR _9861_ (
    .CLK(clk_bF$buf106),
    .D(_663_[18]),
    .Q(\datapath_1.regfile_1.regOut[11] [18]),
    .R(rst_bF$buf0),
    .S(vdd)
);

OR2X2 _9441_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_519_)
);

OR2X2 _9021_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_299_)
);

NOR3X1 _12498_ (
    .A(\control_1.reg_state.dout [1]),
    .B(\control_1.reg_state.dout [2]),
    .C(\control_1.reg_state.dout [3]),
    .Y(ALUSrcB[0])
);

OR2X2 _12078_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_1857_)
);

FILL FILL_1__14161_ (
);

OR2X2 _18724_ (
    .A(_7627_),
    .B(_7628_),
    .Y(_7629_)
);

FILL FILL_0__18439_ (
);

OR2X2 _18304_ (
    .A(_7215_),
    .B(_7214_),
    .Y(_7216_)
);

FILL FILL_0__18019_ (
);

FILL FILL_0__13154_ (
);

FILL FILL248520x44460 (
);

FILL FILL432440x44460 (
);

FILL FILL_0__9901_ (
);

FILL FILL_1__15786_ (
);

OR2X2 _19509_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8375_)
);

AND2X2 _14644_ (
    .A(_3815_),
    .B(_3814_),
    .Y(_3804_[5])
);

OR2X2 _14224_ (
    .A(MemToReg_bF$buf4),
    .B(ALUOut[27]),
    .Y(_3594_)
);

FILL FILL79800x365560 (
);

FILL FILL466640x266760 (
);

FILL FILL_0__15720_ (
);

FILL FILL_0__15300_ (
);

FILL FILL_0__18192_ (
);

FILL FILL297160x167960 (
);

AND2X2 _15849_ (
    .A(_4225__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_4798_)
);

FILL FILL155800x306280 (
);

AND2X2 _15429_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_4384_)
);

FILL FILL384560x172900 (
);

DFFSR _15009_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[28]),
    .Q(\datapath_1.PCJump [28]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL312360x212420 (
);

OR2X2 _10984_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .B(_1322__bF$buf3),
    .Y(_1308_)
);

FILL FILL_0__10699_ (
);

OR2X2 _10564_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_1124__bF$buf0),
    .Y(_1088_)
);

FILL FILL_0__10279_ (
);

OR2X2 _10144_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_926__bF$buf1),
    .Y(_868_)
);

FILL FILL_0__16925_ (
);

FILL FILL_0__16505_ (
);

FILL FILL_0__11640_ (
);

FILL FILL323760x281580 (
);

FILL FILL_0__19397_ (
);

AND2X2 _19262_ (
    .A(_6300__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_8159_)
);

DFFSR _8712_ (
    .CLK(clk_bF$buf32),
    .D(_69_[30]),
    .Q(\datapath_1.regfile_1.regOut[2] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL_1__18717_ (
);

OR2X2 _11769_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_1711_)
);

OR2X2 _11349_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_1491_)
);

FILL FILL91200x133380 (
);

FILL FILL_0__12845_ (
);

OR2X2 _12710_ (
    .A(_2269_),
    .B(_2274_),
    .Y(_2275_)
);

FILL FILL_0__12005_ (
);

FILL FILL291080x242060 (
);

OR2X2 _15182_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_4140_)
);

AND2X2 _9917_ (
    .A(_756_),
    .B(_755_),
    .Y(_729_[13])
);

FILL FILL377720x217360 (
);

FILL FILL458280x54340 (
);

INVX1 _13915_ (
    .A(ALUSrcB[0]),
    .Y(_3346_)
);

FILL FILL278160x113620 (
);

AND2X2 _16387_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_5327_)
);

FILL FILL_1__18470_ (
);

FILL FILL_1__9239_ (
);

FILL FILL_0__17043_ (
);

FILL FILL_1__10557_ (
);

FILL FILL494760x44460 (
);

FILL FILL117040x316160 (
);

OR2X2 _9670_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .B(_662__bF$buf4),
    .Y(_632_)
);

OR2X2 _9250_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .B(_464__bF$buf2),
    .Y(_412_)
);

FILL FILL103360x340860 (
);

FILL FILL_0__18668_ (
);

OR2X2 _18953_ (
    .A(_7853_),
    .B(_7854_),
    .Y(_7855_)
);

FILL FILL_0__18248_ (
);

AND2X2 _18533_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_7441_)
);

OR2X2 _18113_ (
    .A(_7027_),
    .B(_7024_),
    .Y(_7028_)
);

FILL FILL_0__13383_ (
);

FILL FILL_1__12703_ (
);

FILL FILL_0__9710_ (
);

FILL FILL_1__15175_ (
);

AND2X2 _19318_ (
    .A(_6272__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_8214_)
);

DFFSR _14873_ (
    .CLK(clk_bF$buf38),
    .D(_3870_[21]),
    .Q(_2_[21]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL_0__14588_ (
);

FILL FILL_0__14168_ (
);

OR2X2 _14453_ (
    .A(vdd),
    .B(\datapath_1.Data [28]),
    .Y(_3728_)
);

AND2X2 _14033_ (
    .A(_3350__bF$buf0),
    .B(_2_[16]),
    .Y(_3448_)
);

FILL FILL259160x4940 (
);

FILL FILL342000x276640 (
);

FILL FILL269800x326040 (
);

AND2X2 _15658_ (
    .A(_4189__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_4610_)
);

AND2X2 _15238_ (
    .A(_4195__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [0]),
    .Y(_4196_)
);

AND2X2 _10793_ (
    .A(_1200_),
    .B(_1199_),
    .Y(_1191_[4])
);

DFFSR _10373_ (
    .CLK(clk_bF$buf21),
    .D(_927_[14]),
    .Q(\datapath_1.regfile_1.regOut[15] [14]),
    .R(rst_bF$buf90),
    .S(vdd)
);

FILL FILL_1__17321_ (
);

FILL FILL_0__10088_ (
);

FILL FILL_0__16314_ (
);

FILL FILL255360x256880 (
);

OR2X2 _19491_ (
    .A(gnd),
    .B(_8385__bF$buf2),
    .Y(_8363_)
);

AND2X2 _19071_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_7971_)
);

FILL FILL443080x148200 (
);

DFFSR _8941_ (
    .CLK(clk_bF$buf85),
    .D(_201_[1]),
    .Q(\datapath_1.regfile_1.regOut[4] [1]),
    .R(rst_bF$buf71),
    .S(vdd)
);

OR2X2 _8521_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_68__bF$buf1),
    .Y(_46_)
);

OR2X2 _11998_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_1850__bF$buf1),
    .Y(_1824_)
);

FILL FILL_1__18946_ (
);

OR2X2 _11578_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .B(_1652__bF$buf2),
    .Y(_1604_)
);

DFFSR _11158_ (
    .CLK(clk_bF$buf81),
    .D(_1323_[25]),
    .Q(\datapath_1.regfile_1.regOut[21] [25]),
    .R(rst_bF$buf13),
    .S(vdd)
);

FILL FILL_0__17939_ (
);

FILL FILL_0__17519_ (
);

INVX1 _17804_ (
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_6723_)
);

FILL FILL_0__12654_ (
);

FILL FILL59280x88920 (
);

DFFSR _9726_ (
    .CLK(clk_bF$buf113),
    .D(_597_[12]),
    .Q(\datapath_1.regfile_1.regOut[10] [12]),
    .R(rst_bF$buf102),
    .S(vdd)
);

OR2X2 _9306_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_449_)
);

FILL FILL203680x59280 (
);

FILL FILL_1__14026_ (
);

AND2X2 _13724_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[19]),
    .Y(_3200_)
);

FILL FILL_0__13019_ (
);

AND2X2 _13304_ (
    .A(_2845_),
    .B(_2843_),
    .Y(_2846_)
);

FILL FILL334400x291460 (
);

OR2X2 _16196_ (
    .A(_5137_),
    .B(_5138_),
    .Y(_5139_)
);

FILL FILL_0__14800_ (
);

FILL FILL431680x242060 (
);

FILL FILL_0__17692_ (
);

FILL FILL_0__17272_ (
);

FILL FILL285760x64220 (
);

AND2X2 _14929_ (
    .A(_3965_),
    .B(_3964_),
    .Y(_3936_[14])
);

AND2X2 _14509_ (
    .A(_3745_),
    .B(_3744_),
    .Y(_3738_[3])
);

FILL FILL53200x330980 (
);

FILL FILL_0__10720_ (
);

FILL FILL_0__10300_ (
);

FILL FILL147440x365560 (
);

FILL FILL_0__18897_ (
);

OR2X2 _18762_ (
    .A(_7665_),
    .B(_7666_),
    .Y(_7667_)
);

FILL FILL_0__18477_ (
);

AND2X2 _18342_ (
    .A(_6321__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_7253_)
);

FILL FILL34200x167960 (
);

FILL FILL348840x118560 (
);

FILL FILL_0__8998_ (
);

OR2X2 _10849_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .B(_1256__bF$buf3),
    .Y(_1238_)
);

OR2X2 _10429_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .B(_1058__bF$buf2),
    .Y(_1018_)
);

OR2X2 _10009_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .B(_860__bF$buf2),
    .Y(_798_)
);

DFFSR _19547_ (
    .CLK(clk_bF$buf6),
    .D(_8320_[24]),
    .Q(\datapath_1.regfile_1.regOut[0] [24]),
    .R(rst_bF$buf34),
    .S(vdd)
);

OR2X2 _19127_ (
    .A(_8025_),
    .B(_8022_),
    .Y(_8026_)
);

OR2X2 _14682_ (
    .A(\datapath_1.rd1 [18]),
    .B(_3869__bF$buf2),
    .Y(_3841_)
);

FILL FILL_0__14397_ (
);

OR2X2 _14262_ (
    .A(\datapath_1.ALUResult [7]),
    .B(_3671__bF$buf3),
    .Y(_3621_)
);

FILL FILL105640x227240 (
);

OR2X2 _15887_ (
    .A(_4834_),
    .B(_4833_),
    .Y(_4835_)
);

OR2X2 _15467_ (
    .A(_4421_),
    .B(_4420_),
    .Y(_4422_)
);

AND2X2 _15047_ (
    .A(_4034_),
    .B(_4035_),
    .Y(_4036_)
);

FILL FILL211280x301340 (
);

FILL FILL_1__17970_ (
);

OR2X2 _10182_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_893_)
);

FILL FILL_0__16963_ (
);

FILL FILL_0__16543_ (
);

FILL FILL_0__16123_ (
);

FILL FILL128440x311220 (
);

FILL FILL386840x286520 (
);

AND2X2 _8750_ (
    .A(_158_),
    .B(_157_),
    .Y(_135_[11])
);

FILL FILL_1__18335_ (
);

AND2X2 _11387_ (
    .A(_1516_),
    .B(_1515_),
    .Y(_1455_[30])
);

FILL FILL_1__13050_ (
);

AND2X2 _17613_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_6535_)
);

FILL FILL_0__12883_ (
);

FILL FILL_0__12463_ (
);

OR2X2 _9955_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .B(_794__bF$buf3),
    .Y(_782_)
);

OR2X2 _9535_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .B(_596__bF$buf3),
    .Y(_562_)
);

OR2X2 _9115_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .B(_398__bF$buf0),
    .Y(_342_)
);

FILL FILL_1__14675_ (
);

AND2X2 _18818_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_7722_)
);

FILL FILL_0_BUFX2_insert351 (
);

FILL FILL_0_BUFX2_insert352 (
);

FILL FILL_0_BUFX2_insert353 (
);

AND2X2 _13953_ (
    .A(_3344__bF$buf3),
    .B(gnd),
    .Y(_3379_)
);

FILL FILL_0_BUFX2_insert354 (
);

FILL FILL_0__13668_ (
);

FILL FILL_0__13248_ (
);

FILL FILL_0_BUFX2_insert355 (
);

AND2X2 _13533_ (
    .A(_3043_),
    .B(_3042_),
    .Y(_1_[14])
);

OR2X2 _13113_ (
    .A(_2665_),
    .B(_2259_),
    .Y(_2666_)
);

FILL FILL_0_BUFX2_insert356 (
);

FILL FILL449920x326040 (
);

FILL FILL_0_BUFX2_insert358 (
);

FILL FILL450680x222300 (
);

FILL FILL_0__17081_ (
);

FILL FILL_1__10175_ (
);

DFFSR _14738_ (
    .CLK(clk_bF$buf41),
    .D(_3804_[15]),
    .Q(\datapath_1.a [15]),
    .R(rst_bF$buf63),
    .S(vdd)
);

OR2X2 _14318_ (
    .A(vdd),
    .B(ALUOut[26]),
    .Y(_3658_)
);

FILL FILL297920x237120 (
);

FILL FILL_0__15814_ (
);

FILL FILL_1__19293_ (
);

AND2X2 _18991_ (
    .A(_6255__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_7892_)
);

FILL FILL_0__18286_ (
);

OR2X2 _18571_ (
    .A(_7477_),
    .B(_7478_),
    .Y(_7479_)
);

OR2X2 _18151_ (
    .A(_7063_),
    .B(_7064_),
    .Y(_7065_)
);

AND2X2 _10658_ (
    .A(_1130_),
    .B(_1129_),
    .Y(_1125_[2])
);

DFFSR _10238_ (
    .CLK(clk_bF$buf25),
    .D(_861_[8]),
    .Q(\datapath_1.regfile_1.regOut[14] [8]),
    .R(rst_bF$buf89),
    .S(vdd)
);

FILL FILL315400x330980 (
);

FILL FILL317680x54340 (
);

OR2X2 _19356_ (
    .A(_8244_),
    .B(_8251_),
    .Y(_8252_)
);

DFFSR _14491_ (
    .CLK(clk_bF$buf23),
    .D(_3672_[26]),
    .Q(\datapath_1.Data [26]),
    .R(rst_bF$buf22),
    .S(vdd)
);

OR2X2 _14071_ (
    .A(_3480_),
    .B(_3477_),
    .Y(\datapath_1.alu_1.ALUInB [21])
);

OR2X2 _8806_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .B(_200__bF$buf3),
    .Y(_196_)
);

FILL FILL_1__13526_ (
);

AND2X2 _12804_ (
    .A(_2363_),
    .B(_2368_),
    .Y(_2369_)
);

FILL FILL_0__12519_ (
);

FILL FILL84360x345800 (
);

FILL FILL345040x192660 (
);

OR2X2 _15696_ (
    .A(_4646_),
    .B(_4643_),
    .Y(_4647_)
);

AND2X2 _15276_ (
    .A(_4207_),
    .B(_4144_),
    .Y(_4234_)
);

FILL FILL255360x326040 (
);

FILL FILL_0__16772_ (
);

FILL FILL_1__18984_ (
);

FILL FILL259160x247000 (
);

OR2X2 _11196_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_1409_)
);

FILL FILL_0__17557_ (
);

AND2X2 _17842_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_6761_)
);

AND2X2 _17422_ (
    .A(_6317__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_6347_)
);

FILL FILL_0__17137_ (
);

AND2X2 _17002_ (
    .A(_4223__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_5933_)
);

FILL FILL_0__12272_ (
);

FILL FILL408120x232180 (
);

AND2X2 _9764_ (
    .A(_674_),
    .B(_673_),
    .Y(_663_[5])
);

DFFSR _9344_ (
    .CLK(clk_bF$buf8),
    .D(_399_[17]),
    .Q(\datapath_1.regfile_1.regOut[7] [17]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL61560x44460 (
);

FILL FILL421800x54340 (
);

AND2X2 _18627_ (
    .A(_6287__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_7534_)
);

AND2X2 _18207_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_7120_)
);

FILL FILL462080x34580 (
);

FILL FILL_0__13897_ (
);

FILL FILL_0__13477_ (
);

AND2X2 _13762_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [24]),
    .Y(_3233_)
);

NOR2X1 _13342_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2882_)
);

FILL FILL214320x54340 (
);

FILL FILL494760x247000 (
);

FILL FILL_0__9804_ (
);

FILL FILL425600x108680 (
);

FILL FILL116280x128440 (
);

OR2X2 _14967_ (
    .A(\datapath_1.mux_pcsrc.dout [27]),
    .B(_4001__bF$buf3),
    .Y(_3991_)
);

FILL FILL321480x306280 (
);

OR2X2 _14547_ (
    .A(memoryOutData[16]),
    .B(_3803__bF$buf4),
    .Y(_3771_)
);

OR2X2 _14127_ (
    .A(_3528_),
    .B(_3525_),
    .Y(\datapath_1.alu_1.ALUInB [29])
);

FILL FILL_0__15623_ (
);

FILL FILL250800x44460 (
);

FILL FILL_0__18095_ (
);

OR2X2 _18380_ (
    .A(_7287_),
    .B(_7290_),
    .Y(_7291_)
);

FILL FILL503880x217360 (
);

FILL FILL41800x14820 (
);

FILL FILL65360x44460 (
);

FILL FILL425600x54340 (
);

FILL FILL237120x167960 (
);

DFFSR _10887_ (
    .CLK(clk_bF$buf113),
    .D(_1191_[12]),
    .Q(\datapath_1.regfile_1.regOut[19] [12]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_1__17835_ (
);

FILL FILL_1__17415_ (
);

OR2X2 _10467_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_1043_)
);

OR2X2 _10047_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_823_)
);

FILL FILL28880x281580 (
);

FILL FILL_0__16408_ (
);

FILL FILL218120x54340 (
);

FILL FILL_0__11963_ (
);

AND2X2 _19165_ (
    .A(_8063_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd1 [27])
);

AND2X2 _8615_ (
    .A(_88_),
    .B(_87_),
    .Y(_69_[9])
);

FILL FILL145160x39520 (
);

FILL FILL290320x256880 (
);

FILL FILL100320x123500 (
);

FILL FILL60040x261820 (
);

FILL FILL_0__12748_ (
);

INVX1 _12613_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2178_)
);

FILL FILL_0__12328_ (
);

FILL FILL374680x212420 (
);

FILL FILL364040x172900 (
);

OR2X2 _15085_ (
    .A(\datapath_1.a3 [4]),
    .B(_4069_),
    .Y(_4070_)
);

FILL FILL45600x14820 (
);

FILL FILL355680x370500 (
);

FILL FILL400520x207480 (
);

FILL FILL_0__16161_ (
);

AND2X2 _13818_ (
    .A(_3278_),
    .B(_3341_),
    .Y(\datapath_1.alu_1.ALUInA [0])
);

FILL FILL_0__17786_ (
);

OR2X2 _17651_ (
    .A(_6565_),
    .B(_6572_),
    .Y(_6573_)
);

FILL FILL_0__17366_ (
);

OR2X2 _17231_ (
    .A(_6156_),
    .B(_6157_),
    .Y(_6158_)
);

FILL FILL440800x301340 (
);

FILL FILL22800x88920 (
);

DFFSR _9993_ (
    .CLK(clk_bF$buf93),
    .D(_729_[21]),
    .Q(\datapath_1.regfile_1.regOut[12] [21]),
    .R(rst_bF$buf38),
    .S(vdd)
);

OR2X2 _9573_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_587_)
);

FILL FILL460560x54340 (
);

OR2X2 _9153_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_367_)
);

FILL FILL_1__19158_ (
);

FILL FILL402800x296400 (
);

AND2X2 _18856_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_7759_)
);

FILL FILL_0_BUFX2_insert731 (
);

AND2X2 _18436_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_7346_)
);

FILL FILL480320x69160 (
);

FILL FILL_0_BUFX2_insert732 (
);

AND2X2 _18016_ (
    .A(_6255__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_6932_)
);

FILL FILL_0_BUFX2_insert733 (
);

AND2X2 _13991_ (
    .A(_3350__bF$buf3),
    .B(_2_[10]),
    .Y(_3412_)
);

FILL FILL_0_BUFX2_insert734 (
);

FILL FILL_0_BUFX2_insert735 (
);

FILL FILL_0__13286_ (
);

OR2X2 _13571_ (
    .A(ALUOut[27]),
    .B(_3079__bF$buf0),
    .Y(_3069_)
);

MUX2X1 _13151_ (
    .A(_2376__bF$buf2),
    .B(_2501_),
    .S(_2458_),
    .Y(_2702_)
);

FILL FILL_0_BUFX2_insert737 (
);

FILL FILL_0_BUFX2_insert739 (
);

FILL FILL44080x24700 (
);

FILL FILL249280x311220 (
);

FILL FILL243200x335920 (
);

AND2X2 _14776_ (
    .A(_3883_),
    .B(_3882_),
    .Y(_3870_[6])
);

DFFSR _14356_ (
    .CLK(clk_bF$buf40),
    .D(_3606_[20]),
    .Q(ALUOut[20]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL_0__15432_ (
);

FILL FILL440800x24700 (
);

FILL FILL186200x286520 (
);

FILL FILL83600x79040 (
);

FILL FILL493240x113620 (
);

OR2X2 _10696_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .B(_1190__bF$buf0),
    .Y(_1156_)
);

OR2X2 _10276_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .B(_992__bF$buf4),
    .Y(_936_)
);

FILL FILL_0__16637_ (
);

AND2X2 _16922_ (
    .A(_4175__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_5854_)
);

OR2X2 _16502_ (
    .A(_5440_),
    .B(_5437_),
    .Y(_5441_)
);

FILL FILL474240x271700 (
);

FILL FILL_0__11772_ (
);

FILL FILL_0__11352_ (
);

FILL FILL402040x311220 (
);

FILL FILL465880x148200 (
);

OR2X2 _19394_ (
    .A(_8287_),
    .B(_8288_),
    .Y(_8289_)
);

INVX2 _8844_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .Y(_266_)
);

BUFX2 _8424_ (
    .A(_2_[0]),
    .Y(memoryWriteData[0])
);

FILL FILL332120x316160 (
);

FILL FILL_1__13564_ (
);

FILL FILL_1__13144_ (
);

OR2X2 _17707_ (
    .A(_6627_),
    .B(_6626_),
    .Y(_6628_)
);

AOI22X1 _12842_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .C(\datapath_1.alu_1.ALUInB [4]),
    .D(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2407_)
);

AND2X2 _12422_ (
    .A(_2046_),
    .B(_2045_),
    .Y(_1983_[31])
);

FILL FILL449160x88920 (
);

AND2X2 _12002_ (
    .A(_1826_),
    .B(_1825_),
    .Y(_1785_[20])
);

FILL FILL25080x98800 (
);

AND2X2 _9629_ (
    .A(_604_),
    .B(_603_),
    .Y(_597_[3])
);

DFFSR _9209_ (
    .CLK(clk_bF$buf79),
    .D(_333_[11]),
    .Q(\datapath_1.regfile_1.regOut[6] [11]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL_0__16390_ (
);

FILL FILL180120x227240 (
);

AND2X2 _13627_ (
    .A(_3084__bF$buf4),
    .B(\aluControl_1.inst [3]),
    .Y(_3117_)
);

NOR2X1 _13207_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2755_)
);

OR2X2 _16099_ (
    .A(_5042_),
    .B(_5043_),
    .Y(_5044_)
);

FILL FILL_0__14703_ (
);

OR2X2 _17880_ (
    .A(_6797_),
    .B(_6794_),
    .Y(_6798_)
);

FILL FILL_0__17595_ (
);

AND2X2 _17460_ (
    .A(_6255__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_6385_)
);

OR2X2 _17040_ (
    .A(_5966_),
    .B(_5969_),
    .Y(_5970_)
);

FILL FILL453720x340860 (
);

FILL FILL81320x311220 (
);

FILL FILL_1__10269_ (
);

OR2X2 _9382_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .B(_530__bF$buf2),
    .Y(_480_)
);

FILL FILL91200x83980 (
);

FILL FILL_1__11630_ (
);

FILL FILL_0__15908_ (
);

FILL FILL_1__19387_ (
);

OR2X2 _18665_ (
    .A(_7568_),
    .B(_7570_),
    .Y(_7571_)
);

AND2X2 _18245_ (
    .A(_6300__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_7158_)
);

FILL FILL440040x345800 (
);

FILL FILL_0__13095_ (
);

AND2X2 _13380_ (
    .A(_2917_),
    .B(_2907_),
    .Y(_2918_)
);

FILL FILL_0__19321_ (
);

FILL FILL_0__9422_ (
);

OR2X2 _14585_ (
    .A(IRWrite_bF$buf2),
    .B(\control_1.op [3]),
    .Y(_3796_)
);

OR2X2 _14165_ (
    .A(\datapath_1.Data [7]),
    .B(_3605__bF$buf0),
    .Y(_3555_)
);

FILL FILL_0__15661_ (
);

FILL FILL_0__15241_ (
);

FILL FILL217360x19760 (
);

FILL FILL_1_BUFX2_insert284 (
);

FILL FILL_1_BUFX2_insert286 (
);

FILL FILL_1_BUFX2_insert288 (
);

FILL FILL41800x217360 (
);

FILL FILL_1__17453_ (
);

AND2X2 _10085_ (
    .A(_848_),
    .B(_847_),
    .Y(_795_[26])
);

FILL FILL309320x276640 (
);

FILL FILL54720x163020 (
);

AND2X2 _16731_ (
    .A(_4200__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_5666_)
);

FILL FILL_0__16026_ (
);

OR2X2 _16311_ (
    .A(_5252_),
    .B(_5245_),
    .Y(_5253_)
);

FILL FILL_0__11581_ (
);

FILL FILL274360x0 (
);

OR2X2 _8653_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .B(_134__bF$buf4),
    .Y(_114_)
);

FILL FILL190000x9880 (
);

FILL FILL290320x326040 (
);

FILL FILL_1__13793_ (
);

OR2X2 _17936_ (
    .A(_6851_),
    .B(_6852_),
    .Y(_6853_)
);

FILL FILL377720x103740 (
);

OR2X2 _17516_ (
    .A(_6438_),
    .B(_6439_),
    .Y(_6440_)
);

FILL FILL_0__12786_ (
);

NAND2X1 _12651_ (
    .A(_2214_),
    .B(_2215_),
    .Y(_2216_)
);

OR2X2 _12231_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_1939_)
);

DFFSR _9858_ (
    .CLK(clk_bF$buf18),
    .D(_663_[15]),
    .Q(\datapath_1.regfile_1.regOut[11] [15]),
    .R(rst_bF$buf107),
    .S(vdd)
);

OR2X2 _9438_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_517_)
);

OR2X2 _9018_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_297_)
);

FILL FILL102600x237120 (
);

OR2X2 _13856_ (
    .A(\datapath_1.a [13]),
    .B(_3342__bF$buf1),
    .Y(_3304_)
);

NAND2X1 _13436_ (
    .A(_2390_),
    .B(_2379__bF$buf2),
    .Y(_2970_)
);

NAND2X1 _13016_ (
    .A(_2547_),
    .B(_2574_),
    .Y(_2575_)
);

FILL FILL_0__14512_ (
);

FILL FILL351120x0 (
);

FILL FILL_1__16304_ (
);

AND2X2 _9191_ (
    .A(_392_),
    .B(_391_),
    .Y(_333_[29])
);

FILL FILL_0__10852_ (
);

FILL FILL_0__10432_ (
);

AND2X2 _18894_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_7797_)
);

OR2X2 _18474_ (
    .A(_7381_),
    .B(_7382_),
    .Y(_7383_)
);

OR2X2 _18054_ (
    .A(_6968_),
    .B(_6969_),
    .Y(_6970_)
);

FILL FILL324520x148200 (
);

FILL FILL_1__17929_ (
);

FILL FILL438520x217360 (
);

FILL FILL_1__12644_ (
);

FILL FILL_0__9651_ (
);

FILL FILL_0__11637_ (
);

FILL FILL_0__9231_ (
);

DFFSR _11922_ (
    .CLK(clk_bF$buf89),
    .D(_1719_[15]),
    .Q(\datapath_1.regfile_1.regOut[27] [15]),
    .R(rst_bF$buf24),
    .S(vdd)
);

OR2X2 _11502_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_1573_)
);

FILL FILL_0__11217_ (
);

OR2X2 _19259_ (
    .A(_8155_),
    .B(_8147_),
    .Y(_8156_)
);

FILL FILL116280x14820 (
);

OR2X2 _14394_ (
    .A(memoryOutData[8]),
    .B(_3737__bF$buf4),
    .Y(_3689_)
);

FILL FILL146680x247000 (
);

DFFSR _8709_ (
    .CLK(clk_bF$buf68),
    .D(_69_[27]),
    .Q(\datapath_1.regfile_1.regOut[2] [27]),
    .R(rst_bF$buf21),
    .S(vdd)
);

FILL FILL_0__15890_ (
);

FILL FILL487160x242060 (
);

FILL FILL_1__13009_ (
);

FILL FILL367840x192660 (
);

INVX1 _12707_ (
    .A(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2272_)
);

OR2X2 _15599_ (
    .A(_4548_),
    .B(_4551_),
    .Y(_4552_)
);

OR2X2 _15179_ (
    .A(_4131_),
    .B(_4136_),
    .Y(_4137_)
);

FILL FILL_0__16675_ (
);

OR2X2 _16960_ (
    .A(_5889_),
    .B(_5890_),
    .Y(_5891_)
);

OR2X2 _16540_ (
    .A(_5477_),
    .B(_5476_),
    .Y(_5478_)
);

FILL FILL_0__16255_ (
);

FILL FILL126160x133380 (
);

OR2X2 _16120_ (
    .A(_5049_),
    .B(_5064_),
    .Y(_5065_)
);

FILL FILL_0__11390_ (
);

FILL FILL459040x375440 (
);

AND2X2 _8882_ (
    .A(_226_),
    .B(_225_),
    .Y(_201_[12])
);

AND2X2 _8462_ (
    .A(_6_),
    .B(_5_),
    .Y(_3_[1])
);

FILL FILL_1__10710_ (
);

AND2X2 _11099_ (
    .A(_1364_),
    .B(_1363_),
    .Y(_1323_[20])
);

FILL FILL108680x306280 (
);

OR2X2 _17745_ (
    .A(_6663_),
    .B(_6664_),
    .Y(_6665_)
);

AND2X2 _17325_ (
    .A(_6250__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_6251_)
);

FILL FILL_0__12595_ (
);

NAND3X1 _12880_ (
    .A(_2417_),
    .B(\datapath_1.alu_1.ALUInB [14]),
    .C(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2445_)
);

INVX1 _12460_ (
    .A(ALUOp[0]),
    .Y(_2054_)
);

DFFSR _12040_ (
    .CLK(clk_bF$buf24),
    .D(_1785_[4]),
    .Q(\datapath_1.regfile_1.regOut[28] [4]),
    .R(rst_bF$buf82),
    .S(vdd)
);

FILL FILL_0__18821_ (
);

FILL FILL_0__18401_ (
);

OR2X2 _9667_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .B(_662__bF$buf4),
    .Y(_630_)
);

OR2X2 _9247_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .B(_464__bF$buf2),
    .Y(_410_)
);

FILL FILL_0__8922_ (
);

FILL FILL_0__10908_ (
);

FILL FILL_0__8502_ (
);

FILL FILL_1_BUFX2_insert1044 (
);

AND2X2 _13665_ (
    .A(_3089__bF$buf4),
    .B(gnd),
    .Y(_3150_)
);

XOR2X1 _13245_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2790_)
);

FILL FILL_1_BUFX2_insert1046 (
);

FILL FILL_1_BUFX2_insert1048 (
);

FILL FILL18240x64220 (
);

FILL FILL316160x256880 (
);

FILL FILL_0__9707_ (
);

FILL FILL284240x311220 (
);

FILL FILL_1__16953_ (
);

FILL FILL_1__16533_ (
);

FILL FILL_0__15526_ (
);

AND2X2 _15811_ (
    .A(_4154__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_4760_)
);

FILL FILL_0__15106_ (
);

FILL FILL_0__10661_ (
);

FILL FILL356440x350740 (
);

OR2X2 _18283_ (
    .A(_7190_),
    .B(_7194_),
    .Y(_7195_)
);

FILL FILL365560x79040 (
);

FILL FILL_0__9040_ (
);

FILL FILL_0__11446_ (
);

OR2X2 _11731_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_1718__bF$buf1),
    .Y(_1686_)
);

FILL FILL338200x83980 (
);

OR2X2 _11311_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .B(_1520__bF$buf2),
    .Y(_1466_)
);

OR2X2 _19488_ (
    .A(gnd),
    .B(_8385__bF$buf4),
    .Y(_8361_)
);

AND2X2 _19068_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_7968_)
);

FILL FILL4560x261820 (
);

OR2X2 _8938_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .B(_266__bF$buf0),
    .Y(_264_)
);

OR2X2 _8518_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .B(_68__bF$buf2),
    .Y(_44_)
);

FILL FILL10640x301340 (
);

FILL FILL_1__13658_ (
);

FILL FILL299440x167960 (
);

FILL FILL227240x207480 (
);

FILL FILL386840x172900 (
);

INVX1 _12936_ (
    .A(ALUControl[1]),
    .Y(_2500_)
);

INVX1 _12516_ (
    .A(_2096_),
    .Y(_2107_)
);

FILL FILL_1_BUFX2_insert664 (
);

FILL FILL_1_BUFX2_insert666 (
);

FILL FILL_1_BUFX2_insert668 (
);

FILL FILL340480x153140 (
);

FILL FILL_0__16484_ (
);

FILL FILL_0__16064_ (
);

FILL FILL257640x163020 (
);

DFFSR _8691_ (
    .CLK(clk_bF$buf113),
    .D(_69_[9]),
    .Q(\datapath_1.regfile_1.regOut[2] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

FILL FILL254600x0 (
);

FILL FILL138320x49400 (
);

FILL FILL130720x335920 (
);

FILL FILL_1__18276_ (
);

BUFX2 BUFX2_insert330 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf1 )
);

BUFX2 BUFX2_insert331 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf0 )
);

BUFX2 BUFX2_insert332 (
    .A(_596_),
    .Y(_596__bF$buf4)
);

BUFX2 BUFX2_insert333 (
    .A(_596_),
    .Y(_596__bF$buf3)
);

BUFX2 BUFX2_insert334 (
    .A(_596_),
    .Y(_596__bF$buf2)
);

OR2X2 _17974_ (
    .A(_6887_),
    .B(_6890_),
    .Y(_6891_)
);

FILL FILL293360x242060 (
);

BUFX2 BUFX2_insert335 (
    .A(_596_),
    .Y(_596__bF$buf1)
);

OR2X2 _17554_ (
    .A(_6473_),
    .B(_6476_),
    .Y(_6477_)
);

BUFX2 BUFX2_insert336 (
    .A(_596_),
    .Y(_596__bF$buf0)
);

OR2X2 _17134_ (
    .A(_6061_),
    .B(_6062_),
    .Y(_6063_)
);

BUFX2 BUFX2_insert337 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf4 )
);

BUFX2 BUFX2_insert338 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf3 )
);

BUFX2 BUFX2_insert339 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf2 )
);

AND2X2 _9896_ (
    .A(_742_),
    .B(_741_),
    .Y(_729_[6])
);

DFFSR _9476_ (
    .CLK(clk_bF$buf57),
    .D(_465_[20]),
    .Q(\datapath_1.regfile_1.regOut[8] [20]),
    .R(rst_bF$buf81),
    .S(vdd)
);

AND2X2 _9056_ (
    .A(_322_),
    .B(_321_),
    .Y(_267_[27])
);

FILL FILL452200x167960 (
);

FILL FILL_0__8731_ (
);

FILL FILL_0__10717_ (
);

FILL FILL504640x335920 (
);

OR2X2 _18759_ (
    .A(_7662_),
    .B(_7663_),
    .Y(_7664_)
);

AND2X2 _18339_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [15]),
    .Y(_7250_)
);

OR2X2 _13894_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [26]),
    .Y(_3329_)
);

FILL FILL63080x113620 (
);

FILL FILL_0__13189_ (
);

OR2X2 _13474_ (
    .A(\datapath_1.PCJump [13]),
    .B(_3005_),
    .Y(_3006_)
);

OAI21X1 _13054_ (
    .A(_2266_),
    .B(_2376__bF$buf2),
    .C(_2610_),
    .Y(_2611_)
);

FILL FILL_0__19415_ (
);

FILL FILL_0__14970_ (
);

FILL FILL_0__14550_ (
);

FILL FILL_0__14130_ (
);

FILL FILL209000x182780 (
);

FILL FILL_0__9936_ (
);

FILL FILL_0__9516_ (
);

FILL FILL119320x316160 (
);

OR2X2 _14679_ (
    .A(\datapath_1.rd1 [17]),
    .B(_3869__bF$buf3),
    .Y(_3839_)
);

OR2X2 _14259_ (
    .A(\datapath_1.ALUResult [6]),
    .B(_3671__bF$buf0),
    .Y(_3619_)
);

FILL FILL105640x340860 (
);

FILL FILL_0__15755_ (
);

OR2X2 _15620_ (
    .A(_4571_),
    .B(_4570_),
    .Y(_4572_)
);

AND2X2 _15200_ (
    .A(_4157_),
    .B(_4144_),
    .Y(_4158_)
);

FILL FILL_0__10470_ (
);

FILL FILL131480x281580 (
);

AND2X2 _18092_ (
    .A(_6259__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_7007_)
);

FILL FILL433200x113620 (
);

FILL FILL232560x4940 (
);

OR2X2 _10599_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_1111_)
);

OR2X2 _10179_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_891_)
);

FILL FILL_1__12682_ (
);

OR2X2 _16825_ (
    .A(_5727_),
    .B(_5758_),
    .Y(_5759_)
);

AND2X2 _16405_ (
    .A(_4172__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_5345_)
);

FILL FILL240920x247000 (
);

FILL FILL57000x49400 (
);

AND2X2 _11960_ (
    .A(_1798_),
    .B(_1797_),
    .Y(_1785_[6])
);

DFFSR _11540_ (
    .CLK(clk_bF$buf9),
    .D(_1521_[20]),
    .Q(\datapath_1.regfile_1.regOut[24] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

AND2X2 _11120_ (
    .A(_1378_),
    .B(_1377_),
    .Y(_1323_[27])
);

AND2X2 _19297_ (
    .A(_6328__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_8193_)
);

FILL FILL_0__17901_ (
);

AND2X2 _8747_ (
    .A(_156_),
    .B(_155_),
    .Y(_135_[10])
);

FILL FILL73720x24700 (
);

NAND2X1 _12745_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(_2261_),
    .Y(_2310_)
);

DFFSR _12325_ (
    .CLK(clk_bF$buf100),
    .D(_1917_[31]),
    .Q(\datapath_1.regfile_1.regOut[30] [31]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL_0__13401_ (
);

FILL FILL257640x256880 (
);

FILL FILL270560x4940 (
);

FILL FILL_1__9430_ (
);

FILL FILL481840x321100 (
);

FILL FILL267520x88920 (
);

FILL FILL451440x88920 (
);

FILL FILL_0__17498_ (
);

AND2X2 _17783_ (
    .A(_6287__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_6703_)
);

FILL FILL_0__17078_ (
);

AND2X2 _17363_ (
    .A(_6235_),
    .B(_6201_),
    .Y(_6289_)
);

FILL FILL202920x29640 (
);

FILL FILL_1__16818_ (
);

OR2X2 _9285_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_435_)
);

FILL FILL17480x29640 (
);

FILL FILL215840x118560 (
);

FILL FILL_0__8540_ (
);

FILL FILL_0__10526_ (
);

AND2X2 _10811_ (
    .A(_1212_),
    .B(_1211_),
    .Y(_1191_[10])
);

AND2X2 _18988_ (
    .A(_6321__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_7889_)
);

OR2X2 _18568_ (
    .A(_7472_),
    .B(_7475_),
    .Y(_7476_)
);

OR2X2 _18148_ (
    .A(_7060_),
    .B(_7061_),
    .Y(_7062_)
);

FILL FILL410400x256880 (
);

NAND3X1 _13283_ (
    .A(_2379__bF$buf1),
    .B(\datapath_1.alu_1.ALUInB [9]),
    .C(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2826_)
);

FILL FILL_0__19224_ (
);

FILL FILL_0__9325_ (
);

DFFSR _14488_ (
    .CLK(clk_bF$buf11),
    .D(_3672_[23]),
    .Q(\datapath_1.Data [23]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _14068_ (
    .A(_3350__bF$buf2),
    .B(_2_[21]),
    .Y(_3478_)
);

FILL FILL450680x158080 (
);

FILL FILL_0__15984_ (
);

FILL FILL_0__15144_ (
);

FILL FILL150480x261820 (
);

FILL FILL_1__12491_ (
);

FILL FILL_0__16769_ (
);

AND2X2 _16634_ (
    .A(_5570_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.rd2 [21])
);

FILL FILL_0__16349_ (
);

OR2X2 _16214_ (
    .A(_5156_),
    .B(_5155_),
    .Y(_5157_)
);

FILL FILL_0__11484_ (
);

FILL FILL214320x9880 (
);

FILL FILL103360x44460 (
);

FILL FILL330600x59280 (
);

FILL FILL95000x330980 (
);

OR2X2 _8976_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_269_)
);

DFFSR _8556_ (
    .CLK(clk_bF$buf45),
    .D(_3_[3]),
    .Q(\datapath_1.regfile_1.regOut[1] [3]),
    .R(rst_bF$buf57),
    .S(vdd)
);

FILL FILL123120x59280 (
);

FILL FILL505400x69160 (
);

AND2X2 _17839_ (
    .A(_6236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_6758_)
);

FILL FILL412680x39520 (
);

AND2X2 _17419_ (
    .A(_6315__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [1]),
    .Y(_6344_)
);

OR2X2 _12974_ (
    .A(_2387__bF$buf1),
    .B(_2535_),
    .Y(_2536_)
);

FILL FILL_0__12689_ (
);

FILL FILL213560x301340 (
);

OR2X2 _12554_ (
    .A(_2140_),
    .B(_2141_),
    .Y(_2142_)
);

AND2X2 _12134_ (
    .A(_1894_),
    .B(_1893_),
    .Y(_1851_[21])
);

FILL FILL233320x9880 (
);

FILL FILL_0__18915_ (
);

FILL FILL_0__13630_ (
);

AND2X2 _13759_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[24]),
    .Y(_3230_)
);

XOR2X1 _13339_ (
    .A(_2848_),
    .B(_2861_),
    .Y(_2879_)
);

FILL FILL_1__15422_ (
);

FILL FILL_0__14835_ (
);

OR2X2 _14700_ (
    .A(\datapath_1.rd1 [24]),
    .B(_3869__bF$buf0),
    .Y(_3853_)
);

FILL FILL_0__14415_ (
);

BUFX2 BUFX2_insert710 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf3 )
);

BUFX2 BUFX2_insert711 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf2 )
);

BUFX2 BUFX2_insert712 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf1 )
);

BUFX2 BUFX2_insert713 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf0 )
);

FILL FILL357200x103740 (
);

BUFX2 BUFX2_insert714 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf4 )
);

BUFX2 BUFX2_insert715 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf3 )
);

OR2X2 _17592_ (
    .A(_6514_),
    .B(_6513_),
    .Y(_6515_)
);

BUFX2 BUFX2_insert716 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf2 )
);

AND2X2 _17172_ (
    .A(_4187__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_6100_)
);

BUFX2 BUFX2_insert717 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf1 )
);

BUFX2 BUFX2_insert718 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf0 )
);

FILL FILL15960x49400 (
);

BUFX2 BUFX2_insert719 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf4 )
);

FILL FILL15200x187720 (
);

FILL FILL503880x330980 (
);

FILL FILL338200x261820 (
);

FILL FILL351120x256880 (
);

DFFSR _9094_ (
    .CLK(clk_bF$buf80),
    .D(_267_[25]),
    .Q(\datapath_1.regfile_1.regOut[5] [25]),
    .R(rst_bF$buf76),
    .S(vdd)
);

FILL FILL_1__11762_ (
);

AND2X2 _15905_ (
    .A(_4217__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_4853_)
);

DFFSR _10620_ (
    .CLK(clk_bF$buf27),
    .D(_1059_[3]),
    .Q(\datapath_1.regfile_1.regOut[17] [3]),
    .R(rst_bF$buf28),
    .S(vdd)
);

OR2X2 _10200_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_905_)
);

AND2X2 _18797_ (
    .A(_6317__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_7701_)
);

AND2X2 _18377_ (
    .A(_6247__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_7288_)
);

OR2X2 _13092_ (
    .A(_2274_),
    .B(_2601_),
    .Y(_2647_)
);

FILL FILL446880x281580 (
);

FILL FILL_0__19033_ (
);

FILL FILL15960x172900 (
);

FILL FILL_1__12127_ (
);

FILL FILL391400x350740 (
);

FILL FILL_0__9554_ (
);

AND2X2 _11825_ (
    .A(_1728_),
    .B(_1727_),
    .Y(_1719_[4])
);

DFFSR _11405_ (
    .CLK(clk_bF$buf63),
    .D(_1455_[14]),
    .Q(\datapath_1.regfile_1.regOut[23] [14]),
    .R(rst_bF$buf60),
    .S(vdd)
);

OR2X2 _14297_ (
    .A(vdd),
    .B(ALUOut[19]),
    .Y(_3644_)
);

FILL FILL_0__12901_ (
);

FILL FILL_0__15793_ (
);

FILL FILL_0__15373_ (
);

FILL FILL_1__8510_ (
);

FILL FILL185440x59280 (
);

FILL FILL_0__16998_ (
);

FILL FILL_0__16578_ (
);

OR2X2 _16863_ (
    .A(_5795_),
    .B(_5794_),
    .Y(_5796_)
);

AND2X2 _16443_ (
    .A(_4130__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_5382_)
);

OR2X2 _16023_ (
    .A(_4968_),
    .B(_4965_),
    .Y(_4969_)
);

FILL FILL262200x207480 (
);

FILL FILL232560x83980 (
);

OR2X2 _8785_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .B(_200__bF$buf2),
    .Y(_182_)
);

FILL FILL8360x345800 (
);

FILL FILL340480x316160 (
);

FILL FILL_1__13085_ (
);

FILL FILL86640x345800 (
);

AND2X2 _17648_ (
    .A(_6264__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_6570_)
);

OR2X2 _17228_ (
    .A(_6153_),
    .B(_6154_),
    .Y(_6155_)
);

AND2X2 _12783_ (
    .A(_2345_),
    .B(_2347_),
    .Y(_2348_)
);

FILL FILL_0__12498_ (
);

FILL FILL_0__12078_ (
);

OR2X2 _12363_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_2007_)
);

FILL FILL_0__18304_ (
);

FILL FILL412680x355680 (
);

FILL FILL_1__11818_ (
);

FILL FILL_0__8405_ (
);

FILL FILL169480x291460 (
);

AND2X2 _13988_ (
    .A(_3344__bF$buf0),
    .B(gnd),
    .Y(_3409_)
);

OR2X2 _13568_ (
    .A(ALUOut[26]),
    .B(_3079__bF$buf4),
    .Y(_3067_)
);

AND2X2 _13148_ (
    .A(_2698_),
    .B(_2697_),
    .Y(_2699_)
);

FILL FILL88920x0 (
);

FILL FILL_1__15651_ (
);

FILL FILL_0__19509_ (
);

FILL FILL367080x321100 (
);

FILL FILL_0__14644_ (
);

FILL FILL_0__14224_ (
);

FILL FILL_1__11571_ (
);

FILL FILL205200x148200 (
);

FILL FILL_0__15849_ (
);

AND2X2 _15714_ (
    .A(_4195__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_4665_)
);

FILL FILL_0__10984_ (
);

FILL FILL20520x64220 (
);

FILL FILL341240x133380 (
);

FILL FILL104120x167960 (
);

OR2X2 _18186_ (
    .A(_7099_),
    .B(_7091_),
    .Y(_7100_)
);

FILL FILL378480x256880 (
);

FILL FILL140600x340860 (
);

FILL FILL_0__19262_ (
);

FILL FILL_1__12776_ (
);

OR2X2 _16919_ (
    .A(_5847_),
    .B(_5850_),
    .Y(_5851_)
);

FILL FILL_0__9783_ (
);

FILL FILL_0__9363_ (
);

FILL FILL_0__11769_ (
);

FILL FILL_0__11349_ (
);

OR2X2 _11634_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_1641_)
);

OR2X2 _11214_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_1421_)
);

FILL FILL_0__12710_ (
);

FILL FILL180880x14820 (
);

FILL FILL_0__15182_ (
);

FILL FILL64600x14820 (
);

FILL FILL281200x321100 (
);

FILL FILL239400x167960 (
);

OR2X2 _12839_ (
    .A(_2401_),
    .B(_2403_),
    .Y(_2404_)
);

AND2X2 _12419_ (
    .A(_2044_),
    .B(_2043_),
    .Y(_1983_[30])
);

FILL FILL72200x316160 (
);

FILL FILL222680x370500 (
);

FILL FILL41040x14820 (
);

FILL FILL_1__17394_ (
);

FILL FILL180880x108680 (
);

OR2X2 _16672_ (
    .A(_5604_),
    .B(_5607_),
    .Y(_5608_)
);

AND2X2 _16252_ (
    .A(_4160__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_5194_)
);

FILL FILL298680x232180 (
);

FILL FILL448400x266760 (
);

FILL FILL210520x158080 (
);

AND2X2 _8594_ (
    .A(_74_),
    .B(_73_),
    .Y(_69_[2])
);

FILL FILL41800x88920 (
);

FILL FILL292600x256880 (
);

FILL FILL_1__10842_ (
);

FILL FILL17480x286520 (
);

FILL FILL62320x261820 (
);

FILL FILL376960x212420 (
);

AND2X2 _17877_ (
    .A(_6326__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_6795_)
);

AND2X2 _17457_ (
    .A(_6259__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_6382_)
);

AND2X2 _17037_ (
    .A(_4230__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_5967_)
);

FILL FILL366320x172900 (
);

OR2X2 _12592_ (
    .A(_2153_),
    .B(_2156_),
    .Y(_2157_)
);

FILL FILL68400x14820 (
);

DFFSR _12172_ (
    .CLK(clk_bF$buf39),
    .D(_1851_[7]),
    .Q(\datapath_1.regfile_1.regOut[29] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

FILL FILL357960x370500 (
);

FILL FILL231800x74100 (
);

FILL FILL_0__18953_ (
);

FILL FILL_0__18533_ (
);

FILL FILL402800x207480 (
);

FILL FILL_0__18113_ (
);

OR2X2 _9799_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .B(_728__bF$buf0),
    .Y(_698_)
);

OR2X2 _9379_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_530__bF$buf2),
    .Y(_478_)
);

FILL FILL431680x335920 (
);

FILL FILL_1__11207_ (
);

FILL FILL_0__8634_ (
);

DFFSR _10905_ (
    .CLK(clk_bF$buf32),
    .D(_1191_[30]),
    .Q(\datapath_1.regfile_1.regOut[19] [30]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL_1__14099_ (
);

FILL FILL116280x311220 (
);

AND2X2 _13797_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [29]),
    .Y(_3263_)
);

XOR2X1 _13377_ (
    .A(_2190_),
    .B(_2400_),
    .Y(_2915_)
);

FILL FILL_1__15040_ (
);

FILL FILL302480x326040 (
);

FILL FILL_0__14033_ (
);

FILL FILL_0__9839_ (
);

FILL FILL28880x143260 (
);

FILL FILL235600x74100 (
);

OR2X2 _15943_ (
    .A(_4888_),
    .B(_4889_),
    .Y(_4890_)
);

FILL FILL_0__15658_ (
);

OR2X2 _15523_ (
    .A(_4475_),
    .B(_4476_),
    .Y(_4477_)
);

FILL FILL_0__15238_ (
);

AND2X2 _15103_ (
    .A(_4041_),
    .B(_4084_),
    .Y(_4085_)
);

FILL FILL_0__10793_ (
);

FILL FILL254600x360620 (
);

FILL FILL_0__19491_ (
);

OR2X2 _16728_ (
    .A(_5655_),
    .B(_5662_),
    .Y(_5663_)
);

AND2X2 _16308_ (
    .A(_4183__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_5250_)
);

FILL FILL_1__18811_ (
);

FILL FILL_0__11578_ (
);

FILL FILL_0__9172_ (
);

OR2X2 _11863_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .B(_1784__bF$buf2),
    .Y(_1754_)
);

OR2X2 _11443_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .B(_1586__bF$buf1),
    .Y(_1534_)
);

DFFSR _11023_ (
    .CLK(clk_bF$buf16),
    .D(_1257_[19]),
    .Q(\datapath_1.regfile_1.regOut[20] [19]),
    .R(rst_bF$buf20),
    .S(vdd)
);

FILL FILL_0__17804_ (
);

FILL FILL85120x355680 (
);

NAND2X1 _12648_ (
    .A(_2211_),
    .B(_2212_),
    .Y(_2213_)
);

OR2X2 _12228_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_1937_)
);

FILL FILL_0__13724_ (
);

FILL FILL404320x311220 (
);

FILL FILL_0_BUFX2_insert1050 (
);

FILL FILL_0_BUFX2_insert1051 (
);

FILL FILL_0_BUFX2_insert1052 (
);

FILL FILL_0_BUFX2_insert1053 (
);

AND2X2 _16481_ (
    .A(_4230__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_5420_)
);

FILL FILL_0__16196_ (
);

OR2X2 _16061_ (
    .A(_5005_),
    .B(_5004_),
    .Y(_5006_)
);

FILL FILL_0_BUFX2_insert1054 (
);

FILL FILL_0_BUFX2_insert1056 (
);

FILL FILL_0_BUFX2_insert1058 (
);

FILL FILL334400x316160 (
);

FILL FILL_1__15516_ (
);

FILL FILL_0__14929_ (
);

FILL FILL389880x251940 (
);

FILL FILL270560x74100 (
);

FILL FILL502360x291460 (
);

FILL FILL246240x281580 (
);

OR2X2 _17686_ (
    .A(_6598_),
    .B(_6606_),
    .Y(_6607_)
);

OR2X2 _17266_ (
    .A(_6191_),
    .B(_6192_),
    .Y(_6193_)
);

FILL FILL252320x222300 (
);

FILL FILL_0__18762_ (
);

FILL FILL_0__18342_ (
);

AND2X2 _9188_ (
    .A(_390_),
    .B(_389_),
    .Y(_333_[28])
);

FILL FILL182400x227240 (
);

FILL FILL382280x0 (
);

FILL FILL_0__8863_ (
);

FILL FILL_0__8443_ (
);

OR2X2 _10714_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_1190__bF$buf3),
    .Y(_1168_)
);

FILL FILL_0__10429_ (
);

FILL FILL_0__10009_ (
);

FILL FILL66120x301340 (
);

XOR2X1 _13186_ (
    .A(_2211_),
    .B(_2734_),
    .Y(_2735_)
);

OR2X2 _19412_ (
    .A(_8305_),
    .B(_8306_),
    .Y(_8307_)
);

FILL FILL_0__19127_ (
);

FILL FILL_0__14682_ (
);

FILL FILL_0__9648_ (
);

DFFSR _11919_ (
    .CLK(clk_bF$buf106),
    .D(_1719_[12]),
    .Q(\datapath_1.regfile_1.regOut[27] [12]),
    .R(rst_bF$buf0),
    .S(vdd)
);

FILL FILL291080x24700 (
);

FILL FILL420280x19760 (
);

FILL FILL_1__16474_ (
);

FILL FILL47880x123500 (
);

OR2X2 _15752_ (
    .A(_4698_),
    .B(_4701_),
    .Y(_4702_)
);

FILL FILL_0__15467_ (
);

FILL FILL_0__15047_ (
);

AND2X2 _15332_ (
    .A(_4154__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_4289_)
);

FILL FILL_0__10182_ (
);

FILL FILL186200x335920 (
);

FILL FILL291840x98800 (
);

FILL FILL_1__17259_ (
);

OR2X2 _16957_ (
    .A(_5887_),
    .B(_5886_),
    .Y(_5888_)
);

OR2X2 _16537_ (
    .A(_5474_),
    .B(_5459_),
    .Y(_5475_)
);

OR2X2 _16117_ (
    .A(_5061_),
    .B(_5060_),
    .Y(_5062_)
);

DFFSR _11672_ (
    .CLK(clk_bF$buf83),
    .D(_1587_[23]),
    .Q(\datapath_1.regfile_1.regOut[25] [23]),
    .R(rst_bF$buf17),
    .S(vdd)
);

AND2X2 _11252_ (
    .A(_1446_),
    .B(_1445_),
    .Y(_1389_[28])
);

FILL FILL_0__17613_ (
);

AND2X2 _8879_ (
    .A(_224_),
    .B(_223_),
    .Y(_201_[11])
);

AND2X2 _8459_ (
    .A(_4_),
    .B(_67_),
    .Y(_3_[0])
);

FILL FILL216600x370500 (
);

OR2X2 _9820_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .B(_728__bF$buf0),
    .Y(_712_)
);

OR2X2 _9400_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .B(_530__bF$buf0),
    .Y(_492_)
);

FILL FILL_1__13599_ (
);

AOI22X1 _12877_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .C(\datapath_1.alu_1.ALUInB [12]),
    .D(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2442_)
);

FILL FILL174800x108680 (
);

AND2X2 _12457_ (
    .A(_2050_),
    .B(\aluControl_1.inst [5]),
    .Y(_2051_)
);

DFFSR _12037_ (
    .CLK(clk_bF$buf43),
    .D(_1785_[1]),
    .Q(\datapath_1.regfile_1.regOut[28] [1]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL_0__18818_ (
);

FILL FILL_0__13533_ (
);

FILL FILL_0__13113_ (
);

FILL FILL295640x98800 (
);

FILL FILL462080x133380 (
);

AND2X2 _16290_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_5232_)
);

FILL FILL_1__9562_ (
);

FILL FILL_1__10460_ (
);

FILL FILL_0__14318_ (
);

DFFSR _14603_ (
    .CLK(clk_bF$buf31),
    .D(_3738_[9]),
    .Q(\datapath_1.PCJump [11]),
    .R(rst_bF$buf85),
    .S(vdd)
);

OR2X2 _17495_ (
    .A(_6417_),
    .B(_6418_),
    .Y(_6419_)
);

AND2X2 _17075_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_6005_)
);

FILL FILL256880x138320 (
);

FILL FILL_0__18991_ (
);

OR2X2 _15808_ (
    .A(_4755_),
    .B(_4756_),
    .Y(_4757_)
);

AND2X2 _10943_ (
    .A(_1280_),
    .B(_1279_),
    .Y(_1257_[11])
);

AND2X2 _10523_ (
    .A(_1060_),
    .B(_1123_),
    .Y(_1059_[0])
);

DFFSR _10103_ (
    .CLK(clk_bF$buf112),
    .D(_795_[2]),
    .Q(\datapath_1.regfile_1.regOut[13] [2]),
    .R(rst_bF$buf3),
    .S(vdd)
);

FILL FILL11400x54340 (
);

FILL FILL9880x227240 (
);

FILL FILL_0__19356_ (
);

FILL FILL118560x64220 (
);

OR2X2 _19221_ (
    .A(_8117_),
    .B(_8118_),
    .Y(_8119_)
);

FILL FILL_0__14071_ (
);

FILL FILL_0__9877_ (
);

FILL FILL217360x182780 (
);

OR2X2 _11728_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .B(_1718__bF$buf0),
    .Y(_1684_)
);

OR2X2 _11308_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .B(_1520__bF$buf4),
    .Y(_1464_)
);

AND2X2 _15981_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_4928_)
);

FILL FILL_0__15696_ (
);

OR2X2 _15561_ (
    .A(_4506_),
    .B(_4513_),
    .Y(_4514_)
);

AND2X2 _15141_ (
    .A(_4109_),
    .B(_4016_),
    .Y(\datapath_1.regfile_1.regEn [21])
);

FILL FILL329840x64220 (
);

FILL FILL237880x0 (
);

FILL FILL_1__17488_ (
);

FILL FILL326040x375440 (
);

AND2X2 _16766_ (
    .A(_4187__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_5700_)
);

AND2X2 _16346_ (
    .A(_4181__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_5287_)
);

OR2X2 _11481_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_1559_)
);

OR2X2 _11061_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_1339_)
);

FILL FILL_0__17422_ (
);

FILL FILL452960x182780 (
);

FILL FILL_0__17002_ (
);

DFFSR _8688_ (
    .CLK(clk_bF$buf32),
    .D(_69_[6]),
    .Q(\datapath_1.regfile_1.regOut[2] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

OR2X2 _12686_ (
    .A(_2250_),
    .B(_2213_),
    .Y(_2251_)
);

AND2X2 _12266_ (
    .A(_1962_),
    .B(_1961_),
    .Y(_1917_[22])
);

FILL FILL_0__18627_ (
);

OR2X2 _18912_ (
    .A(_7810_),
    .B(_7813_),
    .Y(_7814_)
);

FILL FILL_0__18207_ (
);

FILL FILL128440x133380 (
);

FILL FILL_0__13762_ (
);

FILL FILL_0__13342_ (
);

FILL FILL178600x69160 (
);

FILL FILL_1__9371_ (
);

FILL FILL505400x182780 (
);

FILL FILL_0__14967_ (
);

OR2X2 _14832_ (
    .A(\datapath_1.rd2 [25]),
    .B(_3935__bF$buf3),
    .Y(_3921_)
);

FILL FILL_0__14547_ (
);

OR2X2 _14412_ (
    .A(memoryOutData[14]),
    .B(_3737__bF$buf3),
    .Y(_3701_)
);

FILL FILL200640x266760 (
);

FILL FILL237120x326040 (
);

FILL FILL_0__18380_ (
);

FILL FILL_1__16339_ (
);

FILL FILL_1__11894_ (
);

OR2X2 _15617_ (
    .A(_4565_),
    .B(_4568_),
    .Y(_4569_)
);

FILL FILL_0__8481_ (
);

FILL FILL_0__10467_ (
);

DFFSR _10752_ (
    .CLK(clk_bF$buf68),
    .D(_1125_[6]),
    .Q(\datapath_1.regfile_1.regOut[18] [6]),
    .R(rst_bF$buf40),
    .S(vdd)
);

FILL FILL_1__17700_ (
);

FILL FILL_0__10047_ (
);

OR2X2 _10332_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_973_)
);

OR2X2 _18089_ (
    .A(_7003_),
    .B(_6996_),
    .Y(_7004_)
);

AND2X2 _19450_ (
    .A(_8335_),
    .B(_8334_),
    .Y(_8320_[7])
);

FILL FILL490200x153140 (
);

OR2X2 _19030_ (
    .A(_7927_),
    .B(_7930_),
    .Y(_7931_)
);

AND2X2 _8900_ (
    .A(_238_),
    .B(_237_),
    .Y(_201_[18])
);

FILL FILL_1__12259_ (
);

FILL FILL_0__9686_ (
);

AND2X2 _11957_ (
    .A(_1796_),
    .B(_1795_),
    .Y(_1785_[5])
);

DFFSR _11537_ (
    .CLK(clk_bF$buf76),
    .D(_1521_[17]),
    .Q(\datapath_1.regfile_1.regOut[24] [17]),
    .R(rst_bF$buf112),
    .S(vdd)
);

AND2X2 _11117_ (
    .A(_1376_),
    .B(_1375_),
    .Y(_1323_[26])
);

FILL FILL_0__12613_ (
);

FILL FILL_1__16092_ (
);

FILL FILL35720x276640 (
);

FILL FILL358720x350740 (
);

OR2X2 _15790_ (
    .A(_4738_),
    .B(_4739_),
    .Y(_4740_)
);

FILL FILL_0__15085_ (
);

AND2X2 _15370_ (
    .A(_4228__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_4326_)
);

FILL FILL_1__14405_ (
);

FILL FILL_0__13818_ (
);

FILL FILL67640x251940 (
);

OR2X2 _16995_ (
    .A(_5925_),
    .B(_5924_),
    .Y(_5926_)
);

AND2X2 _16575_ (
    .A(_4130__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_5512_)
);

AND2X2 _16155_ (
    .A(_4200__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_5099_)
);

FILL FILL6840x261820 (
);

DFFSR _11290_ (
    .CLK(clk_bF$buf25),
    .D(_1389_[28]),
    .Q(\datapath_1.regfile_1.regOut[22] [28]),
    .R(rst_bF$buf55),
    .S(vdd)
);

FILL FILL_0__17651_ (
);

FILL FILL_0__17231_ (
);

FILL FILL12920x301340 (
);

OR2X2 _8497_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_68__bF$buf1),
    .Y(_30_)
);

FILL FILL6080x167960 (
);

FILL FILL316920x212420 (
);

FILL FILL12160x207480 (
);

NAND2X1 _12495_ (
    .A(\control_1.reg_state.dout [2]),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2097_)
);

FILL FILL_1__19023_ (
);

OR2X2 _12075_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_1855_)
);

FILL FILL342760x153140 (
);

FILL FILL_0__18856_ (
);

OR2X2 _18721_ (
    .A(_7625_),
    .B(_7624_),
    .Y(_7626_)
);

OR2X2 _18301_ (
    .A(_7205_),
    .B(_7212_),
    .Y(_7213_)
);

FILL FILL_0__13991_ (
);

FILL FILL_0__13571_ (
);

FILL FILL_0__13151_ (
);

FILL FILL281200x281580 (
);

FILL FILL_0__8537_ (
);

FILL FILL278160x232180 (
);

FILL FILL414960x192660 (
);

AND2X2 _10808_ (
    .A(_1210_),
    .B(_1209_),
    .Y(_1191_[9])
);

FILL FILL_1__9180_ (
);

OR2X2 _19506_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8373_)
);

FILL FILL295640x242060 (
);

FILL FILL_0__14776_ (
);

AND2X2 _14641_ (
    .A(_3813_),
    .B(_3812_),
    .Y(_3804_[4])
);

OR2X2 _14221_ (
    .A(MemToReg_bF$buf3),
    .B(ALUOut[26]),
    .Y(_3592_)
);

FILL FILL164160x350740 (
);

FILL FILL337440x370500 (
);

FILL FILL_1__16988_ (
);

OR2X2 _15846_ (
    .A(_4794_),
    .B(_4793_),
    .Y(_4795_)
);

AND2X2 _15426_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_4381_)
);

DFFSR _15006_ (
    .CLK(clk_bF$buf12),
    .D(_3936_[25]),
    .Q(\datapath_1.mux_iord.din0 [25]),
    .R(rst_bF$buf5),
    .S(vdd)
);

OR2X2 _10981_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .B(_1322__bF$buf3),
    .Y(_1306_)
);

OR2X2 _10561_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .B(_1124__bF$buf0),
    .Y(_1086_)
);

FILL FILL_0__10276_ (
);

OR2X2 _10141_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .B(_926__bF$buf1),
    .Y(_866_)
);

FILL FILL300200x113620 (
);

FILL FILL_0__16922_ (
);

FILL FILL_0__16502_ (
);

FILL FILL_0__19394_ (
);

FILL FILL449920x286520 (
);

FILL FILL_1__12068_ (
);

FILL FILL363280x177840 (
);

FILL FILL299440x350740 (
);

FILL FILL221920x316160 (
);

FILL FILL_0__9495_ (
);

OR2X2 _11766_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_1709_)
);

OR2X2 _11346_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_1489_)
);

FILL FILL_0__17707_ (
);

FILL FILL_0__12842_ (
);

FILL FILL_0__12422_ (
);

FILL FILL_0__12002_ (
);

FILL FILL421040x4940 (
);

FILL FILL386080x261820 (
);

AND2X2 _9914_ (
    .A(_754_),
    .B(_753_),
    .Y(_729_[12])
);

FILL FILL_1__8871_ (
);

FILL FILL_1__14214_ (
);

INVX1 _13912_ (
    .A(ALUSrcB[1]),
    .Y(_3343_)
);

FILL FILL_0__13207_ (
);

FILL FILL_0__16099_ (
);

OR2X2 _16384_ (
    .A(_5322_),
    .B(_5323_),
    .Y(_5324_)
);

FILL FILL_0__17880_ (
);

FILL FILL_0__17460_ (
);

FILL FILL40280x212420 (
);

FILL FILL_1__15839_ (
);

FILL FILL65360x4940 (
);

FILL FILL344280x123500 (
);

BUFX2 BUFX2_insert680 (
    .A(_4189_),
    .Y(_4189__bF$buf4)
);

BUFX2 BUFX2_insert681 (
    .A(_4189_),
    .Y(_4189__bF$buf3)
);

BUFX2 BUFX2_insert682 (
    .A(_4189_),
    .Y(_4189__bF$buf2)
);

FILL FILL51680x281580 (
);

BUFX2 BUFX2_insert683 (
    .A(_4189_),
    .Y(_4189__bF$buf1)
);

BUFX2 BUFX2_insert684 (
    .A(_4189_),
    .Y(_4189__bF$buf0)
);

OR2X2 _17589_ (
    .A(_6510_),
    .B(_6511_),
    .Y(_6512_)
);

BUFX2 BUFX2_insert685 (
    .A(_4210_),
    .Y(_4210__bF$buf4)
);

BUFX2 BUFX2_insert686 (
    .A(_4210_),
    .Y(_4210__bF$buf3)
);

AND2X2 _17169_ (
    .A(_4181__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_6097_)
);

BUFX2 BUFX2_insert687 (
    .A(_4210_),
    .Y(_4210__bF$buf2)
);

BUFX2 BUFX2_insert688 (
    .A(_4210_),
    .Y(_4210__bF$buf1)
);

BUFX2 BUFX2_insert689 (
    .A(_4210_),
    .Y(_4210__bF$buf0)
);

FILL FILL_1__19252_ (
);

OR2X2 _18950_ (
    .A(_7844_),
    .B(_7851_),
    .Y(_7852_)
);

FILL FILL_0__18245_ (
);

OR2X2 _18530_ (
    .A(_7433_),
    .B(_7437_),
    .Y(_7438_)
);

AND2X2 _18110_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_7025_)
);

FILL FILL_0__8766_ (
);

DFFSR _10617_ (
    .CLK(clk_bF$buf19),
    .D(_1059_[0]),
    .Q(\datapath_1.regfile_1.regOut[17] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

NAND3X1 _13089_ (
    .A(_2155_),
    .B(ALUControl[0]),
    .C(_2153_),
    .Y(_2644_)
);

FILL FILL_1__15592_ (
);

OR2X2 _19315_ (
    .A(_8209_),
    .B(_8210_),
    .Y(_8211_)
);

FILL FILL452960x0 (
);

DFFSR _14870_ (
    .CLK(clk_bF$buf98),
    .D(_3870_[18]),
    .Q(_2_[18]),
    .R(rst_bF$buf87),
    .S(vdd)
);

FILL FILL_0__14165_ (
);

OR2X2 _14450_ (
    .A(vdd),
    .B(\datapath_1.Data [27]),
    .Y(_3726_)
);

AND2X2 _14030_ (
    .A(_3344__bF$buf2),
    .B(gnd),
    .Y(_3445_)
);

FILL FILL269040x345800 (
);

FILL FILL_1__13905_ (
);

OR2X2 _15655_ (
    .A(_4606_),
    .B(_4603_),
    .Y(_4607_)
);

OR2X2 _15235_ (
    .A(_4192_),
    .B(_4180_),
    .Y(_4193_)
);

AND2X2 _10790_ (
    .A(_1198_),
    .B(_1197_),
    .Y(_1191_[3])
);

DFFSR _10370_ (
    .CLK(clk_bF$buf46),
    .D(_927_[11]),
    .Q(\datapath_1.regfile_1.regOut[15] [11]),
    .R(rst_bF$buf97),
    .S(vdd)
);

FILL FILL249280x133380 (
);

FILL FILL_0__16731_ (
);

FILL FILL504640x54340 (
);

OR2X2 _11995_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .B(_1850__bF$buf4),
    .Y(_1822_)
);

OR2X2 _11575_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .B(_1652__bF$buf1),
    .Y(_1602_)
);

FILL FILL_1__18103_ (
);

DFFSR _11155_ (
    .CLK(clk_bF$buf101),
    .D(_1323_[22]),
    .Q(\datapath_1.regfile_1.regOut[21] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

FILL FILL171760x103740 (
);

FILL FILL229520x29640 (
);

FILL FILL_0__17936_ (
);

AND2X2 _17801_ (
    .A(_6323__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_6720_)
);

FILL FILL_0__12651_ (
);

FILL FILL_0__12231_ (
);

FILL FILL152760x261820 (
);

DFFSR _9723_ (
    .CLK(clk_bF$buf89),
    .D(_597_[9]),
    .Q(\datapath_1.regfile_1.regOut[10] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

OR2X2 _9303_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_447_)
);

FILL FILL344280x350740 (
);

FILL FILL_0__13856_ (
);

FILL FILL_0__13436_ (
);

AND2X2 _13721_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3198_)
);

AND2X2 _13301_ (
    .A(_2842_),
    .B(_2840_),
    .Y(_2843_)
);

FILL FILL_0__13016_ (
);

FILL FILL15200x232180 (
);

FILL FILL402040x133380 (
);

FILL FILL102600x14820 (
);

OR2X2 _16193_ (
    .A(_5132_),
    .B(_5135_),
    .Y(_5136_)
);

FILL FILL34960x49400 (
);

FILL FILL435480x39520 (
);

AND2X2 _14926_ (
    .A(_3963_),
    .B(_3962_),
    .Y(_3936_[13])
);

AND2X2 _14506_ (
    .A(_3743_),
    .B(_3742_),
    .Y(_3738_[2])
);

FILL FILL215840x301340 (
);

FILL FILL461320x9880 (
);

AND2X2 _17398_ (
    .A(_6323__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_6324_)
);

FILL FILL241680x242060 (
);

FILL FILL_0__18894_ (
);

FILL FILL_0__18474_ (
);

FILL FILL_0__18054_ (
);

FILL FILL_0__8995_ (
);

OR2X2 _10846_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .B(_1256__bF$buf3),
    .Y(_1236_)
);

OR2X2 _10426_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_1058__bF$buf0),
    .Y(_1016_)
);

OR2X2 _10006_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_860__bF$buf4),
    .Y(_796_)
);

FILL FILL106400x14820 (
);

FILL FILL_0__11502_ (
);

DFFSR _19544_ (
    .CLK(clk_bF$buf34),
    .D(_8320_[21]),
    .Q(\datapath_1.regfile_1.regOut[0] [21]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_0__19259_ (
);

AND2X2 _19124_ (
    .A(_6262__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_8023_)
);

FILL FILL_0__12707_ (
);

FILL FILL427120x172900 (
);

FILL FILL_0__15599_ (
);

OR2X2 _15884_ (
    .A(_4831_),
    .B(_4830_),
    .Y(_4832_)
);

FILL FILL281960x202540 (
);

OR2X2 _15464_ (
    .A(_4411_),
    .B(_4418_),
    .Y(_4419_)
);

FILL FILL_0__15179_ (
);

NAND3X1 _15044_ (
    .A(_4024_),
    .B(\datapath_1.a3 [4]),
    .C(_4018_),
    .Y(_4033_)
);

FILL FILL_0__16540_ (
);

FILL FILL_0__16120_ (
);

FILL FILL357200x177840 (
);

FILL FILL76000x350740 (
);

FILL FILL198360x118560 (
);

FILL FILL68400x4940 (
);

AND2X2 _16669_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_5605_)
);

OR2X2 _16249_ (
    .A(_5160_),
    .B(_5191_),
    .Y(_5192_)
);

FILL FILL_1__18752_ (
);

FILL FILL426360x93860 (
);

AND2X2 _11384_ (
    .A(_1514_),
    .B(_1513_),
    .Y(_1455_[29])
);

FILL FILL_0__17745_ (
);

AND2X2 _17610_ (
    .A(_6293__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_6532_)
);

FILL FILL_0__17325_ (
);

FILL FILL_0__12880_ (
);

FILL FILL81320x34580 (
);

FILL FILL_0__12460_ (
);

FILL FILL188480x44460 (
);

OR2X2 _9952_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .B(_794__bF$buf2),
    .Y(_780_)
);

OR2X2 _9532_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .B(_596__bF$buf2),
    .Y(_560_)
);

OR2X2 _9112_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .B(_398__bF$buf1),
    .Y(_340_)
);

FILL FILL11400x128440 (
);

INVX1 _12589_ (
    .A(ALUControl[0]),
    .Y(_2154_)
);

DFFSR _12169_ (
    .CLK(clk_bF$buf83),
    .D(_1851_[4]),
    .Q(\datapath_1.regfile_1.regOut[29] [4]),
    .R(rst_bF$buf17),
    .S(vdd)
);

FILL FILL_1__19117_ (
);

AND2X2 _18815_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_7719_)
);

FILL FILL_0_BUFX2_insert321 (
);

FILL FILL_0_BUFX2_insert323 (
);

AND2X2 _13950_ (
    .A(_3352__bF$buf4),
    .B(\aluControl_1.inst [2]),
    .Y(_3377_)
);

FILL FILL_0__13665_ (
);

FILL FILL_0_BUFX2_insert325 (
);

AND2X2 _13530_ (
    .A(_3041_),
    .B(_3040_),
    .Y(_1_[13])
);

AND2X2 _13110_ (
    .A(_2663_),
    .B(_2655_),
    .Y(_2664_)
);

FILL FILL_0_BUFX2_insert327 (
);

FILL FILL_0_BUFX2_insert328 (
);

FILL FILL_0_BUFX2_insert329 (
);

FILL FILL161120x29640 (
);

FILL FILL205960x256880 (
);

FILL FILL_1__9274_ (
);

FILL FILL351120x118560 (
);

FILL FILL_1__15457_ (
);

FILL FILL_1__10592_ (
);

FILL FILL88920x345800 (
);

DFFSR _14735_ (
    .CLK(clk_bF$buf58),
    .D(_3804_[12]),
    .Q(\datapath_1.a [12]),
    .R(rst_bF$buf15),
    .S(vdd)
);

OR2X2 _14315_ (
    .A(vdd),
    .B(ALUOut[25]),
    .Y(_3656_)
);

FILL FILL505400x296400 (
);

FILL FILL500840x98800 (
);

FILL FILL414960x355680 (
);

FILL FILL109440x98800 (
);

AND2X2 _10655_ (
    .A(_1128_),
    .B(_1127_),
    .Y(_1125_[1])
);

DFFSR _10235_ (
    .CLK(clk_bF$buf59),
    .D(_861_[5]),
    .Q(\datapath_1.regfile_1.regOut[14] [5]),
    .R(rst_bF$buf25),
    .S(vdd)
);

FILL FILL285000x365560 (
);

FILL FILL180120x187720 (
);

FILL FILL_0__11731_ (
);

FILL FILL_0__11311_ (
);

FILL FILL_0__19068_ (
);

AND2X2 _19353_ (
    .A(_6236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_8249_)
);

OR2X2 _8803_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .B(_200__bF$buf0),
    .Y(_194_)
);

FILL FILL_0__12936_ (
);

NAND3X1 _12801_ (
    .A(_2365_),
    .B(\datapath_1.alu_1.ALUInA [28]),
    .C(_2364_),
    .Y(_2366_)
);

FILL FILL307040x281580 (
);

FILL FILL43320x64220 (
);

FILL FILL106400x167960 (
);

AND2X2 _15693_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_4644_)
);

AND2X2 _15273_ (
    .A(_4230__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_4231_)
);

FILL FILL_1__8545_ (
);

FILL FILL_1__14308_ (
);

AND2X2 _16898_ (
    .A(_4189__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_5830_)
);

AND2X2 _16478_ (
    .A(_4189__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_5417_)
);

FILL FILL155040x192660 (
);

AND2X2 _16058_ (
    .A(_5003_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd2 [12])
);

FILL FILL_1__18141_ (
);

OR2X2 _11193_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_1407_)
);

FILL FILL_0__17974_ (
);

FILL FILL207480x360620 (
);

FILL FILL_1__10228_ (
);

FILL FILL34960x207480 (
);

AND2X2 _9761_ (
    .A(_672_),
    .B(_671_),
    .Y(_663_[4])
);

DFFSR _9341_ (
    .CLK(clk_bF$buf106),
    .D(_399_[14]),
    .Q(\datapath_1.regfile_1.regOut[7] [14]),
    .R(rst_bF$buf96),
    .S(vdd)
);

AND2X2 _12398_ (
    .A(_2030_),
    .B(_2029_),
    .Y(_1983_[23])
);

FILL FILL_0__18759_ (
);

OR2X2 _18624_ (
    .A(_7529_),
    .B(_7530_),
    .Y(_7531_)
);

FILL FILL_0__18339_ (
);

OR2X2 _18204_ (
    .A(_7116_),
    .B(_7113_),
    .Y(_7117_)
);

FILL FILL_0__13054_ (
);

FILL FILL19760x286520 (
);

FILL FILL64600x261820 (
);

FILL FILL_0__9801_ (
);

OR2X2 _19409_ (
    .A(_8302_),
    .B(_8303_),
    .Y(_8304_)
);

OR2X2 _14964_ (
    .A(\datapath_1.mux_pcsrc.dout [26]),
    .B(_4001__bF$buf1),
    .Y(_3989_)
);

FILL FILL_0__14679_ (
);

FILL FILL368600x172900 (
);

FILL FILL_0__14259_ (
);

OR2X2 _14544_ (
    .A(memoryOutData[15]),
    .B(_3803__bF$buf3),
    .Y(_3769_)
);

FILL FILL41040x88920 (
);

AND2X2 _14124_ (
    .A(_3350__bF$buf2),
    .B(_2_[29]),
    .Y(_3526_)
);

FILL FILL154280x4940 (
);

FILL FILL104120x350740 (
);

FILL FILL_0__15620_ (
);

FILL FILL_0__15200_ (
);

FILL FILL433960x335920 (
);

FILL FILL_0__18092_ (
);

FILL FILL231040x74100 (
);

AND2X2 _15749_ (
    .A(_4234__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_4699_)
);

AND2X2 _15329_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_4286_)
);

FILL FILL131480x306280 (
);

DFFSR _10884_ (
    .CLK(clk_bF$buf55),
    .D(_1191_[9]),
    .Q(\datapath_1.regfile_1.regOut[19] [9]),
    .R(rst_bF$buf27),
    .S(vdd)
);

FILL FILL_0__10599_ (
);

FILL FILL_0__10179_ (
);

OR2X2 _10464_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_1041_)
);

OR2X2 _10044_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_821_)
);

FILL FILL_0__16825_ (
);

FILL FILL_0__16405_ (
);

FILL FILL_0__11120_ (
);

FILL FILL_0__19297_ (
);

OR2X2 _19162_ (
    .A(_8044_),
    .B(_8060_),
    .Y(_8061_)
);

FILL FILL408120x355680 (
);

AND2X2 _8612_ (
    .A(_86_),
    .B(_85_),
    .Y(_69_[8])
);

FILL FILL_0__9398_ (
);

DFFSR _11669_ (
    .CLK(clk_bF$buf27),
    .D(_1587_[20]),
    .Q(\datapath_1.regfile_1.regOut[25] [20]),
    .R(rst_bF$buf28),
    .S(vdd)
);

FILL FILL_1__18617_ (
);

AND2X2 _11249_ (
    .A(_1444_),
    .B(_1443_),
    .Y(_1389_[27])
);

FILL FILL_1__13332_ (
);

FILL FILL13680x227240 (
);

INVX1 _12610_ (
    .A(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2175_)
);

AND2X2 _15082_ (
    .A(_4041_),
    .B(_4067_),
    .Y(_4068_)
);

FILL FILL387600x158080 (
);

OR2X2 _9817_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .B(_728__bF$buf4),
    .Y(_710_)
);

FILL FILL_1__14957_ (
);

OR2X2 _13815_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .B(ALUSrcA_bF$buf0),
    .Y(_3341_)
);

FILL FILL273600x276640 (
);

OR2X2 _16287_ (
    .A(_5227_),
    .B(_5228_),
    .Y(_5229_)
);

FILL FILL_1__18790_ (
);

FILL FILL_1__18370_ (
);

FILL FILL370880x227240 (
);

FILL FILL_0__17363_ (
);

FILL FILL_1__10037_ (
);

DFFSR _9990_ (
    .CLK(clk_bF$buf52),
    .D(_729_[18]),
    .Q(\datapath_1.regfile_1.regOut[12] [18]),
    .R(rst_bF$buf1),
    .S(vdd)
);

OR2X2 _9570_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_585_)
);

OR2X2 _9150_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_365_)
);

FILL FILL478800x271700 (
);

FILL FILL_0__10811_ (
);

FILL FILL406600x311220 (
);

FILL FILL_0__18988_ (
);

FILL FILL_0__18568_ (
);

OR2X2 _18853_ (
    .A(_7754_),
    .B(_7755_),
    .Y(_7756_)
);

FILL FILL_0_BUFX2_insert701 (
);

FILL FILL_0__18148_ (
);

AND2X2 _18433_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_7343_)
);

AND2X2 _18013_ (
    .A(_6321__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_6929_)
);

FILL FILL_0_BUFX2_insert703 (
);

FILL FILL_0_BUFX2_insert705 (
);

FILL FILL_0__13283_ (
);

FILL FILL_0_BUFX2_insert707 (
);

FILL FILL_0_BUFX2_insert708 (
);

FILL FILL_0_BUFX2_insert709 (
);

FILL FILL328320x34580 (
);

FILL FILL_0__8669_ (
);

FILL FILL218880x54340 (
);

FILL FILL256120x98800 (
);

FILL FILL110960x83980 (
);

FILL FILL504640x291460 (
);

FILL FILL_1__15075_ (
);

FILL FILL248520x281580 (
);

OR2X2 _19218_ (
    .A(_8112_),
    .B(_8115_),
    .Y(_8116_)
);

FILL FILL167200x217360 (
);

AND2X2 _14773_ (
    .A(_3881_),
    .B(_3880_),
    .Y(_3870_[5])
);

FILL FILL254600x222300 (
);

DFFSR _14353_ (
    .CLK(clk_bF$buf40),
    .D(_3606_[17]),
    .Q(ALUOut[17]),
    .R(rst_bF$buf53),
    .S(vdd)
);

FILL FILL31160x281580 (
);

FILL FILL74480x345800 (
);

AND2X2 _15978_ (
    .A(_4236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_4925_)
);

AND2X2 _15558_ (
    .A(_4223__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_4511_)
);

NAND2X1 _15138_ (
    .A(_4023_),
    .B(_4043_),
    .Y(_4107_)
);

OR2X2 _10693_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .B(_1190__bF$buf3),
    .Y(_1154_)
);

OR2X2 _10273_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .B(_992__bF$buf0),
    .Y(_934_)
);

FILL FILL_1__17221_ (
);

FILL FILL_0__16214_ (
);

FILL FILL466640x19760 (
);

FILL FILL161880x355680 (
);

AND2X2 _19391_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_8286_)
);

DFFSR _8841_ (
    .CLK(clk_bF$buf7),
    .D(_135_[30]),
    .Q(\datapath_1.regfile_1.regOut[3] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

BUFX2 _8421_ (
    .A(_1_[29]),
    .Y(memoryAddress[29])
);

FILL FILL427120x335920 (
);

FILL FILL259160x19760 (
);

OR2X2 _11898_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_1777_)
);

OR2X2 _11478_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_1557_)
);

OR2X2 _11058_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_1337_)
);

FILL FILL_1__13981_ (
);

FILL FILL_0__17839_ (
);

FILL FILL_0__17419_ (
);

OR2X2 _17704_ (
    .A(_6623_),
    .B(_6624_),
    .Y(_6625_)
);

FILL FILL194560x9880 (
);

FILL FILL_0__12974_ (
);

FILL FILL_0__12554_ (
);

FILL FILL_0__12134_ (
);

AND2X2 _9626_ (
    .A(_602_),
    .B(_601_),
    .Y(_597_[2])
);

DFFSR _9206_ (
    .CLK(clk_bF$buf13),
    .D(_333_[8]),
    .Q(\datapath_1.regfile_1.regOut[6] [8]),
    .R(rst_bF$buf1),
    .S(vdd)
);

FILL FILL_1__14766_ (
);

FILL FILL387600x296400 (
);

AND2X2 _18909_ (
    .A(_6271__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_7811_)
);

FILL FILL291080x98800 (
);

OR2X2 _13624_ (
    .A(_3114_),
    .B(_3113_),
    .Y(_3115_)
);

INVX1 _13204_ (
    .A(_2752_),
    .Y(\datapath_1.ALUResult [15])
);

OR2X2 _16096_ (
    .A(_5037_),
    .B(_5040_),
    .Y(_5041_)
);

FILL FILL_0__17592_ (
);

FILL FILL_0__17172_ (
);

OR2X2 _14829_ (
    .A(\datapath_1.rd2 [24]),
    .B(_3935__bF$buf2),
    .Y(_3919_)
);

OR2X2 _14409_ (
    .A(memoryOutData[13]),
    .B(_3737__bF$buf4),
    .Y(_3699_)
);

FILL FILL_1__16912_ (
);

FILL FILL237880x207480 (
);

FILL FILL_0__15905_ (
);

FILL FILL_0__10200_ (
);

FILL FILL_0__18797_ (
);

AND2X2 _18662_ (
    .A(_6216__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_7568_)
);

FILL FILL_0__18377_ (
);

OR2X2 _18242_ (
    .A(_7154_),
    .B(_7153_),
    .Y(_7155_)
);

FILL FILL_0__13092_ (
);

FILL FILL504640x9880 (
);

FILL FILL_0__8898_ (
);

FILL FILL_0__8478_ (
);

DFFSR _10749_ (
    .CLK(clk_bF$buf27),
    .D(_1125_[3]),
    .Q(\datapath_1.regfile_1.regOut[18] [3]),
    .R(rst_bF$buf28),
    .S(vdd)
);

OR2X2 _10329_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_971_)
);

FILL FILL250040x0 (
);

FILL FILL_1__12412_ (
);

FILL FILL350360x251940 (
);

FILL FILL_0__11825_ (
);

FILL FILL323000x69160 (
);

AND2X2 _19447_ (
    .A(_8333_),
    .B(_8332_),
    .Y(_8320_[6])
);

AND2X2 _19027_ (
    .A(_6302__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_7928_)
);

FILL FILL_0__14297_ (
);

OR2X2 _14582_ (
    .A(IRWrite_bF$buf2),
    .B(\control_1.op [2]),
    .Y(_3794_)
);

OR2X2 _14162_ (
    .A(\datapath_1.Data [6]),
    .B(_3605__bF$buf0),
    .Y(_3553_)
);

FILL FILL280440x256880 (
);

FILL FILL197600x266760 (
);

FILL FILL354160x172900 (
);

FILL FILL_1_BUFX2_insert251 (
);

OR2X2 _15787_ (
    .A(_4736_),
    .B(_4735_),
    .Y(_4737_)
);

OR2X2 _15367_ (
    .A(_4322_),
    .B(_4321_),
    .Y(_4323_)
);

FILL FILL_1__17870_ (
);

AND2X2 _10082_ (
    .A(_846_),
    .B(_845_),
    .Y(_795_[25])
);

FILL FILL275880x375440 (
);

FILL FILL_0__16863_ (
);

FILL FILL_0__16443_ (
);

FILL FILL342000x281580 (
);

FILL FILL180880x335920 (
);

OR2X2 _8650_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .B(_134__bF$buf0),
    .Y(_112_)
);

FILL FILL98040x256880 (
);

FILL FILL_1__18235_ (
);

DFFSR _11287_ (
    .CLK(clk_bF$buf43),
    .D(_1389_[25]),
    .Q(\datapath_1.regfile_1.regOut[22] [25]),
    .R(rst_bF$buf62),
    .S(vdd)
);

OR2X2 _17933_ (
    .A(_6848_),
    .B(_6849_),
    .Y(_6850_)
);

FILL FILL_0__17228_ (
);

OR2X2 _17513_ (
    .A(_6436_),
    .B(_6433_),
    .Y(_6437_)
);

FILL FILL_0__12783_ (
);

FILL FILL_0__12363_ (
);

FILL FILL91960x83980 (
);

DFFSR _9855_ (
    .CLK(clk_bF$buf93),
    .D(_663_[12]),
    .Q(\datapath_1.regfile_1.regOut[11] [12]),
    .R(rst_bF$buf41),
    .S(vdd)
);

OR2X2 _9435_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_515_)
);

OR2X2 _9015_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_295_)
);

OR2X2 _18718_ (
    .A(_7618_),
    .B(_7622_),
    .Y(_7623_)
);

OR2X2 _13853_ (
    .A(\datapath_1.a [12]),
    .B(_3342__bF$buf3),
    .Y(_3302_)
);

FILL FILL_0__13568_ (
);

FILL FILL_0__13148_ (
);

NAND2X1 _13433_ (
    .A(_2853_),
    .B(_2178_),
    .Y(_2967_)
);

OR2X2 _13013_ (
    .A(_2335_),
    .B(_2475_),
    .Y(_2572_)
);

FILL FILL373920x118560 (
);

FILL FILL159600x9880 (
);

FILL FILL73720x128440 (
);

AND2X2 _14638_ (
    .A(_3811_),
    .B(_3810_),
    .Y(_3804_[3])
);

OR2X2 _14218_ (
    .A(MemToReg_bF$buf3),
    .B(ALUOut[25]),
    .Y(_3590_)
);

FILL FILL_0__15714_ (
);

FILL FILL_1__19193_ (
);

FILL FILL483360x113620 (
);

AND2X2 _18891_ (
    .A(_6238__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_7794_)
);

FILL FILL_0__18186_ (
);

OR2X2 _18471_ (
    .A(_7375_),
    .B(_7379_),
    .Y(_7380_)
);

OR2X2 _18051_ (
    .A(_6965_),
    .B(_6966_),
    .Y(_6967_)
);

OR2X2 _10978_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .B(_1322__bF$buf2),
    .Y(_1304_)
);

OR2X2 _10558_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .B(_1124__bF$buf3),
    .Y(_1084_)
);

OR2X2 _10138_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .B(_926__bF$buf2),
    .Y(_864_)
);

FILL FILL_1__12221_ (
);

FILL FILL_0__16919_ (
);

FILL FILL_0__11634_ (
);

AND2X2 _19256_ (
    .A(_6297__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_8153_)
);

FILL FILL202920x266760 (
);

OR2X2 _14391_ (
    .A(memoryOutData[7]),
    .B(_3737__bF$buf4),
    .Y(_3687_)
);

DFFSR _8706_ (
    .CLK(clk_bF$buf97),
    .D(_69_[24]),
    .Q(\datapath_1.regfile_1.regOut[2] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL111720x98800 (
);

FILL FILL_1__13846_ (
);

FILL FILL_1__13426_ (
);

XOR2X1 _12704_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2269_)
);

FILL FILL_0__12419_ (
);

AND2X2 _15596_ (
    .A(_4189__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_4549_)
);

AND2X2 _15176_ (
    .A(_4133_),
    .B(_4128_),
    .Y(_4134_)
);

FILL FILL_0__16672_ (
);

OR2X2 _13909_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.PCJump [31]),
    .Y(_3339_)
);

FILL FILL_1__18884_ (
);

AND2X2 _11096_ (
    .A(_1362_),
    .B(_1361_),
    .Y(_1323_[19])
);

FILL FILL369360x281580 (
);

FILL FILL424840x177840 (
);

FILL FILL_0__17877_ (
);

FILL FILL_0__17457_ (
);

OR2X2 _17742_ (
    .A(_6661_),
    .B(_6658_),
    .Y(_6662_)
);

FILL FILL_0__17037_ (
);

AND2X2 _17322_ (
    .A(_6247__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [0]),
    .Y(_6248_)
);

OR2X2 _9664_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .B(_662__bF$buf1),
    .Y(_628_)
);

OR2X2 _9244_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .B(_464__bF$buf3),
    .Y(_408_)
);

AND2X2 _18947_ (
    .A(_6238__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_7849_)
);

NOR2X1 _18527_ (
    .A(_6310__bF$buf3),
    .B(_7434_),
    .Y(_7435_)
);

AND2X2 _18107_ (
    .A(_6287__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_7022_)
);

FILL FILL_1_BUFX2_insert1011 (
);

FILL FILL_0__13797_ (
);

FILL FILL_0__13377_ (
);

AND2X2 _13662_ (
    .A(_3084__bF$buf3),
    .B(\datapath_1.PCJump [10]),
    .Y(_3147_)
);

AND2X2 _13242_ (
    .A(_2787_),
    .B(_2785_),
    .Y(_2788_)
);

FILL FILL_1_BUFX2_insert1019 (
);

FILL FILL8360x167960 (
);

FILL FILL_0__9704_ (
);

FILL FILL401280x108680 (
);

DFFSR _14867_ (
    .CLK(clk_bF$buf77),
    .D(_3870_[15]),
    .Q(_2_[15]),
    .R(rst_bF$buf65),
    .S(vdd)
);

OR2X2 _14447_ (
    .A(vdd),
    .B(\datapath_1.Data [26]),
    .Y(_3724_)
);

AND2X2 _14027_ (
    .A(_3352__bF$buf0),
    .B(\datapath_1.PCJump [15]),
    .Y(_3443_)
);

FILL FILL_0__15943_ (
);

FILL FILL_0__15523_ (
);

NOR2X1 _18280_ (
    .A(_6310__bF$buf3),
    .B(_7191_),
    .Y(_7192_)
);

FILL FILL_1__11089_ (
);

FILL FILL380760x232180 (
);

AND2X2 _10787_ (
    .A(_1196_),
    .B(_1195_),
    .Y(_1191_[2])
);

FILL FILL_1__17735_ (
);

DFFSR _10367_ (
    .CLK(clk_bF$buf61),
    .D(_927_[8]),
    .Q(\datapath_1.regfile_1.regOut[15] [8]),
    .R(rst_bF$buf58),
    .S(vdd)
);

FILL FILL370120x192660 (
);

FILL FILL316920x286520 (
);

FILL FILL_0__16308_ (
);

FILL FILL_0__11863_ (
);

FILL FILL_0__11443_ (
);

OR2X2 _19485_ (
    .A(gnd),
    .B(_8385__bF$buf1),
    .Y(_8359_)
);

OR2X2 _19065_ (
    .A(_7951_),
    .B(_7964_),
    .Y(_7965_)
);

FILL FILL166440x350740 (
);

OR2X2 _8935_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .B(_266__bF$buf3),
    .Y(_262_)
);

OR2X2 _8515_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .B(_68__bF$buf4),
    .Y(_42_)
);

FILL FILL33440x19760 (
);

FILL FILL288040x64220 (
);

FILL FILL284240x247000 (
);

FILL FILL_1_BUFX2_insert631 (
);

OR2X2 _12933_ (
    .A(_2157__bF$buf0),
    .B(_2496_),
    .Y(_2497_)
);

FILL FILL_0__12648_ (
);

NOR3X1 _12513_ (
    .A(_2102_),
    .B(\control_1.reg_state.dout [2]),
    .C(\control_1.reg_state.dout [3]),
    .Y(_2106_)
);

FILL FILL_0__12228_ (
);

FILL FILL_1_BUFX2_insert639 (
);

FILL FILL_1__8677_ (
);

FILL FILL61560x266760 (
);

FILL FILL_0__16481_ (
);

FILL FILL_0__16061_ (
);

FILL FILL365560x177840 (
);

AND2X2 _13718_ (
    .A(_3084__bF$buf0),
    .B(\datapath_1.PCJump [18]),
    .Y(_3195_)
);

FILL FILL_1__18693_ (
);

BUFX2 BUFX2_insert300 (
    .A(_3737_),
    .Y(_3737__bF$buf2)
);

BUFX2 BUFX2_insert301 (
    .A(_3737_),
    .Y(_3737__bF$buf1)
);

FILL FILL65360x187720 (
);

BUFX2 BUFX2_insert302 (
    .A(_3737_),
    .Y(_3737__bF$buf0)
);

BUFX2 BUFX2_insert303 (
    .A(_332_),
    .Y(_332__bF$buf4)
);

AND2X2 _17971_ (
    .A(_6300__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_6888_)
);

BUFX2 BUFX2_insert304 (
    .A(_332_),
    .Y(_332__bF$buf3)
);

FILL FILL_0__17686_ (
);

FILL FILL_0__17266_ (
);

AND2X2 _17551_ (
    .A(_6271__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_6474_)
);

BUFX2 BUFX2_insert305 (
    .A(_332_),
    .Y(_332__bF$buf2)
);

BUFX2 BUFX2_insert306 (
    .A(_332_),
    .Y(_332__bF$buf1)
);

OR2X2 _17131_ (
    .A(_6058_),
    .B(_6059_),
    .Y(_6060_)
);

BUFX2 BUFX2_insert307 (
    .A(_332_),
    .Y(_332__bF$buf0)
);

BUFX2 BUFX2_insert308 (
    .A(_68_),
    .Y(_68__bF$buf4)
);

BUFX2 BUFX2_insert309 (
    .A(_68_),
    .Y(_68__bF$buf3)
);

FILL FILL300200x187720 (
);

FILL FILL82840x197600 (
);

AND2X2 _9893_ (
    .A(_740_),
    .B(_739_),
    .Y(_729_[5])
);

DFFSR _9473_ (
    .CLK(clk_bF$buf0),
    .D(_465_[17]),
    .Q(\datapath_1.regfile_1.regOut[8] [17]),
    .R(rst_bF$buf64),
    .S(vdd)
);

AND2X2 _9053_ (
    .A(_320_),
    .B(_319_),
    .Y(_267_[26])
);

FILL FILL_1__19058_ (
);

FILL FILL_0__10714_ (
);

OR2X2 _18756_ (
    .A(_7660_),
    .B(_7653_),
    .Y(_7661_)
);

OR2X2 _18336_ (
    .A(_7239_),
    .B(_7246_),
    .Y(_7247_)
);

OR2X2 _13891_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [25]),
    .Y(_3327_)
);

AND2X2 _13471_ (
    .A(_3003_),
    .B(_2982_),
    .Y(ALUZero)
);

NOR2X1 _13051_ (
    .A(_2265_),
    .B(_2498_),
    .Y(_2608_)
);

FILL FILL145160x370500 (
);

FILL FILL_0__9933_ (
);

FILL FILL_0__9513_ (
);

FILL FILL_1__15398_ (
);

OR2X2 _14676_ (
    .A(\datapath_1.rd1 [16]),
    .B(_3869__bF$buf3),
    .Y(_3837_)
);

OR2X2 _14256_ (
    .A(\datapath_1.ALUResult [5]),
    .B(_3671__bF$buf3),
    .Y(_3617_)
);

FILL FILL357960x192660 (
);

FILL FILL_0__15332_ (
);

FILL FILL299440x212420 (
);

FILL FILL84360x0 (
);

OR2X2 _10596_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_1109_)
);

OR2X2 _10176_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_889_)
);

FILL FILL479560x59280 (
);

FILL FILL_0__16957_ (
);

FILL FILL_0__16537_ (
);

OR2X2 _16822_ (
    .A(_5752_),
    .B(_5755_),
    .Y(_5756_)
);

AND2X2 _16402_ (
    .A(_4167__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_5342_)
);

FILL FILL_0__11252_ (
);

OR2X2 _19294_ (
    .A(_8157_),
    .B(_8190_),
    .Y(_8191_)
);

AND2X2 _8744_ (
    .A(_154_),
    .B(_153_),
    .Y(_135_[9])
);

FILL FILL_1__13464_ (
);

AND2X2 _17607_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_6529_)
);

OR2X2 _12742_ (
    .A(_2269_),
    .B(_2306_),
    .Y(_2307_)
);

DFFSR _12322_ (
    .CLK(clk_bF$buf110),
    .D(_1917_[28]),
    .Q(\datapath_1.regfile_1.regOut[30] [28]),
    .R(rst_bF$buf74),
    .S(vdd)
);

OR2X2 _9949_ (
    .A(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .B(_794__bF$buf3),
    .Y(_778_)
);

OR2X2 _9529_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .B(_596__bF$buf0),
    .Y(_558_)
);

OR2X2 _9109_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_398__bF$buf1),
    .Y(_338_)
);

FILL FILL351880x133380 (
);

FILL FILL_0__16290_ (
);

FILL FILL237880x9880 (
);

FILL FILL_0_BUFX2_insert290 (
);

FILL FILL_0_BUFX2_insert291 (
);

FILL FILL_0_BUFX2_insert292 (
);

FILL FILL_0_BUFX2_insert293 (
);

AND2X2 _13947_ (
    .A(_3347__bF$buf0),
    .B(\aluControl_1.inst [4]),
    .Y(_3374_)
);

FILL FILL_0_BUFX2_insert294 (
);

AND2X2 _13527_ (
    .A(_3039_),
    .B(_3038_),
    .Y(_1_[12])
);

XOR2X1 _13107_ (
    .A(_2635_),
    .B(_2615_),
    .Y(_2661_)
);

FILL FILL_0_BUFX2_insert296 (
);

FILL FILL_0_BUFX2_insert298 (
);

FILL FILL329080x340860 (
);

FILL FILL274360x311220 (
);

FILL FILL_0__17495_ (
);

OR2X2 _17780_ (
    .A(_6699_),
    .B(_6696_),
    .Y(_6700_)
);

OR2X2 _17360_ (
    .A(_6284_),
    .B(_6285_),
    .Y(_6286_)
);

FILL FILL256880x9880 (
);

FILL FILL346560x350740 (
);

FILL FILL291840x321100 (
);

OR2X2 _9282_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_433_)
);

FILL FILL_1__11950_ (
);

FILL FILL_1__11110_ (
);

FILL FILL_0__15808_ (
);

FILL FILL_0__10943_ (
);

FILL FILL_0__10523_ (
);

OR2X2 _18985_ (
    .A(_7885_),
    .B(_7878_),
    .Y(_7886_)
);

AND2X2 _18565_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_7473_)
);

OR2X2 _18145_ (
    .A(_7055_),
    .B(_7058_),
    .Y(_7059_)
);

OR2X2 _13280_ (
    .A(_2387__bF$buf3),
    .B(_2822_),
    .Y(_2823_)
);

FILL FILL22800x93860 (
);

FILL FILL_0__19221_ (
);

FILL FILL421800x143260 (
);

FILL FILL112480x163020 (
);

FILL FILL55480x251940 (
);

FILL FILL57760x49400 (
);

FILL FILL458280x39520 (
);

DFFSR _14485_ (
    .CLK(clk_bF$buf78),
    .D(_3672_[20]),
    .Q(\datapath_1.Data [20]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _14065_ (
    .A(_3344__bF$buf4),
    .B(gnd),
    .Y(_3475_)
);

FILL FILL220400x256880 (
);

FILL FILL490960x148200 (
);

FILL FILL243960x242060 (
);

FILL FILL217360x207480 (
);

FILL FILL_0__15561_ (
);

FILL FILL247760x163020 (
);

FILL FILL_1__17353_ (
);

OR2X2 _16631_ (
    .A(_5560_),
    .B(_5567_),
    .Y(_5568_)
);

FILL FILL_0__16346_ (
);

OR2X2 _16211_ (
    .A(_5153_),
    .B(_5152_),
    .Y(_5154_)
);

FILL FILL_0__11481_ (
);

FILL FILL_0__11061_ (
);

FILL FILL_1__9903_ (
);

INVX2 _8973_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .Y(_332_)
);

DFFSR _8553_ (
    .CLK(clk_bF$buf96),
    .D(_3_[0]),
    .Q(\datapath_1.regfile_1.regOut[1] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

FILL FILL38000x256880 (
);

FILL FILL_1__10801_ (
);

FILL FILL_1__18558_ (
);

AND2X2 _17836_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_6755_)
);

OR2X2 _17416_ (
    .A(_6339_),
    .B(_6340_),
    .Y(_6341_)
);

OAI21X1 _12971_ (
    .A(_2357_),
    .B(_2498_),
    .C(_2532_),
    .Y(_2533_)
);

FILL FILL_0__12686_ (
);

FILL FILL_0__12266_ (
);

NOR3X1 _12551_ (
    .A(_2111_),
    .B(\control_1.op [0]),
    .C(_2133_),
    .Y(_2139_)
);

AND2X2 _12131_ (
    .A(_1892_),
    .B(_1891_),
    .Y(_1851_[20])
);

AND2X2 _9758_ (
    .A(_670_),
    .B(_669_),
    .Y(_663_[3])
);

DFFSR _9338_ (
    .CLK(clk_bF$buf95),
    .D(_399_[11]),
    .Q(\datapath_1.regfile_1.regOut[7] [11]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL163400x79040 (
);

FILL FILL465120x251940 (
);

FILL FILL_1__14898_ (
);

AND2X2 _13756_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3228_)
);

FILL FILL144400x153140 (
);

AOI21X1 _13336_ (
    .A(_2547_),
    .B(_2876_),
    .C(_2870_),
    .Y(_2877_)
);

FILL FILL70680x123500 (
);

FILL FILL109440x316160 (
);

FILL FILL505400x207480 (
);

DFFSR _9091_ (
    .CLK(clk_bF$buf26),
    .D(_267_[22]),
    .Q(\datapath_1.regfile_1.regOut[5] [22]),
    .R(rst_bF$buf98),
    .S(vdd)
);

FILL FILL_1__16204_ (
);

AND2X2 _15902_ (
    .A(_4189__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_4850_)
);

FILL FILL_0__10332_ (
);

OR2X2 _18794_ (
    .A(_7696_),
    .B(_7697_),
    .Y(_7698_)
);

AND2X2 _18374_ (
    .A(_6238__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_7285_)
);

FILL FILL_0__19450_ (
);

FILL FILL434720x182780 (
);

FILL FILL_1__12964_ (
);

FILL FILL_1__12544_ (
);

FILL FILL158080x207480 (
);

FILL FILL_0__9971_ (
);

FILL FILL_0__11957_ (
);

AND2X2 _11822_ (
    .A(_1726_),
    .B(_1725_),
    .Y(_1719_[3])
);

FILL FILL_0__9131_ (
);

DFFSR _11402_ (
    .CLK(clk_bF$buf71),
    .D(_1455_[11]),
    .Q(\datapath_1.regfile_1.regOut[23] [11]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL_0__11117_ (
);

OR2X2 _19159_ (
    .A(_8057_),
    .B(_8056_),
    .Y(_8058_)
);

OR2X2 _14294_ (
    .A(vdd),
    .B(ALUOut[18]),
    .Y(_3642_)
);

FILL FILL123880x59280 (
);

AND2X2 _8609_ (
    .A(_84_),
    .B(_83_),
    .Y(_69_[7])
);

FILL FILL_0__15790_ (
);

XOR2X1 _12607_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2172_)
);

FILL FILL182400x187720 (
);

AND2X2 _15499_ (
    .A(_4167__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_4453_)
);

INVX2 _15079_ (
    .A(RegWrite),
    .Y(_4065_)
);

FILL FILL_0__16995_ (
);

OR2X2 _16860_ (
    .A(_5791_),
    .B(_5792_),
    .Y(_5793_)
);

OR2X2 _16440_ (
    .A(_5379_),
    .B(_5364_),
    .Y(_5380_)
);

FILL FILL_0__16155_ (
);

AND2X2 _16020_ (
    .A(_4181__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_4966_)
);

FILL FILL259920x9880 (
);

OR2X2 _8782_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .B(_200__bF$buf1),
    .Y(_180_)
);

FILL FILL11400x311220 (
);

FILL FILL309320x281580 (
);

FILL FILL345800x133380 (
);

AND2X2 _17645_ (
    .A(_6315__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_6567_)
);

OR2X2 _17225_ (
    .A(_6151_),
    .B(_6144_),
    .Y(_6152_)
);

NAND3X1 _12780_ (
    .A(_2325_),
    .B(\datapath_1.alu_1.ALUInA [26]),
    .C(_2344_),
    .Y(_2345_)
);

FILL FILL_0__12495_ (
);

OR2X2 _12360_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_2005_)
);

FILL FILL_0__18721_ (
);

FILL FILL_0__18301_ (
);

DFFSR _9987_ (
    .CLK(clk_bF$buf90),
    .D(_729_[15]),
    .Q(\datapath_1.regfile_1.regOut[12] [15]),
    .R(rst_bF$buf107),
    .S(vdd)
);

OR2X2 _9567_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_583_)
);

OR2X2 _9147_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[6] [15]),
    .Y(_363_)
);

FILL FILL_0__10808_ (
);

FILL FILL_0__8402_ (
);

FILL FILL167960x232180 (
);

FILL FILL_1__14287_ (
);

FILL FILL_0_BUFX2_insert670 (
);

FILL FILL_0_BUFX2_insert671 (
);

FILL FILL_0_BUFX2_insert672 (
);

FILL FILL_0_BUFX2_insert673 (
);

AND2X2 _13985_ (
    .A(_3352__bF$buf0),
    .B(\datapath_1.PCJump [9]),
    .Y(_3407_)
);

FILL FILL_0_BUFX2_insert674 (
);

OR2X2 _13565_ (
    .A(ALUOut[25]),
    .B(_3079__bF$buf1),
    .Y(_3065_)
);

INVX1 _13145_ (
    .A(_2282_),
    .Y(_2696_)
);

FILL FILL_0_BUFX2_insert676 (
);

FILL FILL_0_BUFX2_insert678 (
);

FILL FILL_0__19506_ (
);

FILL FILL60040x88920 (
);

FILL FILL26600x167960 (
);

FILL FILL_1__16853_ (
);

FILL FILL_0__15426_ (
);

OR2X2 _15711_ (
    .A(_4660_),
    .B(_4661_),
    .Y(_4662_)
);

FILL FILL226480x276640 (
);

FILL FILL_0__10561_ (
);

FILL FILL_0__10141_ (
);

AND2X2 _18183_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_7097_)
);

FILL FILL_1__12353_ (
);

AND2X2 _16916_ (
    .A(_4181__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [26]),
    .Y(_5848_)
);

FILL FILL_0__11766_ (
);

OR2X2 _11631_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_1639_)
);

OR2X2 _11211_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_1419_)
);

OR2X2 _19388_ (
    .A(_8282_),
    .B(_8279_),
    .Y(_8283_)
);

FILL FILL106400x350740 (
);

FILL FILL89680x153140 (
);

FILL FILL461320x74100 (
);

DFFSR _8838_ (
    .CLK(clk_bF$buf36),
    .D(_135_[27]),
    .Q(\datapath_1.regfile_1.regOut[3] [27]),
    .R(rst_bF$buf78),
    .S(vdd)
);

BUFX2 _8418_ (
    .A(_1_[26]),
    .Y(memoryAddress[26])
);

FILL FILL188480x256880 (
);

OR2X2 _12836_ (
    .A(_2186_),
    .B(_2187_),
    .Y(_2401_)
);

AND2X2 _12416_ (
    .A(_2042_),
    .B(_2041_),
    .Y(_1983_[29])
);

FILL FILL_0__13912_ (
);

FILL FILL484880x360620 (
);

FILL FILL_0__16384_ (
);

FILL FILL_1__9521_ (
);

FILL FILL235600x59280 (
);

AND2X2 _8591_ (
    .A(_72_),
    .B(_71_),
    .Y(_69_[1])
);

FILL FILL_1__15704_ (
);

FILL FILL_1__18176_ (
);

NOR2X1 _17874_ (
    .A(_6310__bF$buf3),
    .B(_6791_),
    .Y(_6792_)
);

OR2X2 _17454_ (
    .A(_6377_),
    .B(_6378_),
    .Y(_6379_)
);

AND2X2 _17034_ (
    .A(_4167__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_5964_)
);

FILL FILL341240x256880 (
);

FILL FILL_0__18950_ (
);

FILL FILL_0__18110_ (
);

FILL FILL51680x306280 (
);

OR2X2 _9796_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .B(_728__bF$buf2),
    .Y(_696_)
);

OR2X2 _9376_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_530__bF$buf2),
    .Y(_476_)
);

FILL FILL19760x148200 (
);

FILL FILL355680x217360 (
);

FILL FILL_0__8631_ (
);

DFFSR _10902_ (
    .CLK(clk_bF$buf49),
    .D(_1191_[27]),
    .Q(\datapath_1.regfile_1.regOut[19] [27]),
    .R(rst_bF$buf66),
    .S(vdd)
);

OR2X2 _18659_ (
    .A(_7561_),
    .B(_7564_),
    .Y(_7565_)
);

OR2X2 _18239_ (
    .A(_7151_),
    .B(_7149_),
    .Y(_7152_)
);

AND2X2 _13794_ (
    .A(_3081__bF$buf4),
    .B(ALUOut[29]),
    .Y(_3260_)
);

NAND3X1 _13374_ (
    .A(ALUControl[1]),
    .B(\datapath_1.alu_1.ALUInB [4]),
    .C(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2912_)
);

FILL FILL_0__13089_ (
);

FILL FILL_0__19315_ (
);

FILL FILL_0__14450_ (
);

FILL FILL_0__14030_ (
);

FILL FILL362520x187720 (
);

FILL FILL_1__12829_ (
);

CLKBUF1 CLKBUF1_insert220 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert221 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert222 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert223 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf0)
);

FILL FILL_0__9836_ (
);

FILL FILL_0__9416_ (
);

DFFSR _14999_ (
    .CLK(clk_bF$buf40),
    .D(_3936_[18]),
    .Q(\datapath_1.mux_iord.din0 [18]),
    .R(rst_bF$buf65),
    .S(vdd)
);

OR2X2 _14579_ (
    .A(IRWrite_bF$buf2),
    .B(\control_1.op [1]),
    .Y(_3792_)
);

OR2X2 _14159_ (
    .A(\datapath_1.Data [5]),
    .B(_3605__bF$buf1),
    .Y(_3551_)
);

FILL FILL184680x286520 (
);

OR2X2 _15940_ (
    .A(_4885_),
    .B(_4886_),
    .Y(_4887_)
);

FILL FILL_0__15655_ (
);

FILL FILL421800x306280 (
);

OR2X2 _15520_ (
    .A(_4470_),
    .B(_4473_),
    .Y(_4474_)
);

AND2X2 _15100_ (
    .A(_4082_),
    .B(_4076_),
    .Y(_4083_)
);

FILL FILL22040x212420 (
);

DFFSR _10499_ (
    .CLK(clk_bF$buf95),
    .D(_993_[11]),
    .Q(\datapath_1.regfile_1.regOut[16] [11]),
    .R(rst_bF$buf9),
    .S(vdd)
);

FILL FILL_1__17027_ (
);

AND2X2 _10079_ (
    .A(_844_),
    .B(_843_),
    .Y(_795_[24])
);

FILL FILL_1__12162_ (
);

AND2X2 _16725_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_5660_)
);

FILL FILL462080x19760 (
);

AND2X2 _16305_ (
    .A(_4200__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_5247_)
);

FILL FILL_0__11995_ (
);

FILL FILL_0__11575_ (
);

OR2X2 _11860_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_1784__bF$buf2),
    .Y(_1752_)
);

OR2X2 _11440_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .B(_1586__bF$buf1),
    .Y(_1532_)
);

DFFSR _11020_ (
    .CLK(clk_bF$buf11),
    .D(_1257_[16]),
    .Q(\datapath_1.regfile_1.regOut[20] [16]),
    .R(rst_bF$buf111),
    .S(vdd)
);

FILL FILL33440x281580 (
);

FILL FILL420280x182780 (
);

AND2X2 _19197_ (
    .A(_6272__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_8095_)
);

FILL FILL_0__17801_ (
);

OR2X2 _8647_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .B(_134__bF$buf4),
    .Y(_110_)
);

FILL FILL237120x286520 (
);

AND2X2 _12645_ (
    .A(_2193_),
    .B(_2209_),
    .Y(_2210_)
);

OR2X2 _12225_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_1935_)
);

FILL FILL88920x29640 (
);

FILL FILL_0__13301_ (
);

FILL FILL_0_BUFX2_insert1021 (
);

FILL FILL_0_BUFX2_insert1023 (
);

FILL FILL_0_BUFX2_insert1025 (
);

FILL FILL_0_BUFX2_insert1026 (
);

FILL FILL347320x4940 (
);

FILL FILL_0_BUFX2_insert1027 (
);

FILL FILL_0_BUFX2_insert1028 (
);

FILL FILL_0_BUFX2_insert1029 (
);

FILL FILL429400x335920 (
);

FILL FILL_1__15933_ (
);

FILL FILL_0__14506_ (
);

FILL FILL_0__17398_ (
);

AND2X2 _17683_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_6604_)
);

OR2X2 _17263_ (
    .A(_6186_),
    .B(_6189_),
    .Y(_6190_)
);

FILL FILL144400x316160 (
);

FILL FILL231800x321100 (
);

FILL FILL_1__16718_ (
);

AND2X2 _9185_ (
    .A(_388_),
    .B(_387_),
    .Y(_333_[27])
);

FILL FILL_1__11853_ (
);

FILL FILL322240x54340 (
);

FILL FILL_0__10846_ (
);

FILL FILL_0__8440_ (
);

OR2X2 _10711_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .B(_1190__bF$buf2),
    .Y(_1166_)
);

FILL FILL_0__10006_ (
);

NOR2X1 _18888_ (
    .A(_6310__bF$buf1),
    .B(_7790_),
    .Y(_7791_)
);

INVX1 _18468_ (
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_7377_)
);

FILL FILL231040x227240 (
);

OR2X2 _18048_ (
    .A(_6960_),
    .B(_6963_),
    .Y(_6964_)
);

FILL FILL111720x177840 (
);

AND2X2 _13183_ (
    .A(_2731_),
    .B(_2250_),
    .Y(_2732_)
);

FILL FILL_0__19124_ (
);

FILL FILL174800x44460 (
);

FILL FILL_0__9645_ (
);

DFFSR _11916_ (
    .CLK(clk_bF$buf87),
    .D(_1719_[9]),
    .Q(\datapath_1.regfile_1.regOut[27] [9]),
    .R(rst_bF$buf2),
    .S(vdd)
);

FILL FILL504640x340860 (
);

OR2X2 _14388_ (
    .A(memoryOutData[6]),
    .B(_3737__bF$buf1),
    .Y(_3685_)
);

FILL FILL79800x232180 (
);

FILL FILL466640x133380 (
);

FILL FILL349600x54340 (
);

FILL FILL_0__15884_ (
);

FILL FILL_0__15464_ (
);

FILL FILL_0__15044_ (
);

FILL FILL_1__8601_ (
);

FILL FILL352640x251940 (
);

FILL FILL_1__17676_ (
);

FILL FILL66120x237120 (
);

FILL FILL389120x311220 (
);

AND2X2 _16954_ (
    .A(_5885_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd2 [26])
);

OR2X2 _16534_ (
    .A(_5470_),
    .B(_5471_),
    .Y(_5472_)
);

FILL FILL_0__16249_ (
);

OR2X2 _16114_ (
    .A(_5057_),
    .B(_5058_),
    .Y(_5059_)
);

FILL FILL_0__11384_ (
);

FILL FILL282720x256880 (
);

FILL FILL_1__9806_ (
);

FILL FILL470440x148200 (
);

AND2X2 _8876_ (
    .A(_222_),
    .B(_221_),
    .Y(_201_[10])
);

OR2X2 _8456_ (
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .Y(_67_)
);

AND2X2 _17739_ (
    .A(_6326__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_6659_)
);

AND2X2 _17319_ (
    .A(_6244__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [0]),
    .Y(_6245_)
);

FILL FILL_0__12589_ (
);

AND2X2 _12874_ (
    .A(_2434_),
    .B(_2438_),
    .Y(_2439_)
);

DFFSR _12454_ (
    .CLK(clk_bF$buf44),
    .D(_1983_[31]),
    .Q(\datapath_1.regfile_1.regOut[31] [31]),
    .R(rst_bF$buf16),
    .S(vdd)
);

OR2X2 _12034_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .B(_1850__bF$buf3),
    .Y(_1848_)
);

FILL FILL_0__18815_ (
);

FILL FILL_0__13950_ (
);

FILL FILL_0__13530_ (
);

FILL FILL_0__8916_ (
);

OR2X2 _13659_ (
    .A(_3144_),
    .B(_3143_),
    .Y(_3145_)
);

FILL FILL240920x118560 (
);

NOR3X1 _13239_ (
    .A(_2782_),
    .B(_2783_),
    .C(_2784_),
    .Y(_2785_)
);

FILL FILL10640x123500 (
);

FILL FILL_1__15322_ (
);

FILL FILL_0__14315_ (
);

DFFSR _14600_ (
    .CLK(clk_bF$buf31),
    .D(_3738_[6]),
    .Q(\datapath_1.PCJump [8]),
    .R(rst_bF$buf85),
    .S(vdd)
);

FILL FILL184680x0 (
);

AND2X2 _17492_ (
    .A(_6247__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_6416_)
);

AND2X2 _17072_ (
    .A(_4142__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_6002_)
);

FILL FILL153520x24700 (
);

FILL FILL157320x355680 (
);

FILL FILL_1__11242_ (
);

FILL FILL462840x163020 (
);

OR2X2 _15805_ (
    .A(_4753_),
    .B(_4752_),
    .Y(_4754_)
);

FILL FILL_0__10655_ (
);

AND2X2 _10940_ (
    .A(_1278_),
    .B(_1277_),
    .Y(_1257_[10])
);

OR2X2 _10520_ (
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .Y(_1123_)
);

AND2X2 _10100_ (
    .A(_858_),
    .B(_857_),
    .Y(_795_[31])
);

OR2X2 _18697_ (
    .A(_7601_),
    .B(_7602_),
    .Y(_7603_)
);

AND2X2 _18277_ (
    .A(_6317__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_7189_)
);

FILL FILL_0__9034_ (
);

OR2X2 _11725_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .B(_1718__bF$buf2),
    .Y(_1682_)
);

OR2X2 _11305_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .B(_1520__bF$buf4),
    .Y(_1462_)
);

OR2X2 _14197_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[18]),
    .Y(_3576_)
);

FILL FILL_0__12801_ (
);

FILL FILL_1__16280_ (
);

FILL FILL398240x108680 (
);

FILL FILL261440x0 (
);

FILL FILL_0__15273_ (
);

FILL FILL_1__8410_ (
);

FILL FILL79040x276640 (
);

FILL FILL324520x316160 (
);

FILL FILL206720x34580 (
);

FILL FILL_0__16898_ (
);

FILL FILL_0__16478_ (
);

AND2X2 _16763_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_5697_)
);

OR2X2 _16343_ (
    .A(_5283_),
    .B(_5280_),
    .Y(_5284_)
);

FILL FILL_0__11193_ (
);

DFFSR _8685_ (
    .CLK(clk_bF$buf10),
    .D(_69_[3]),
    .Q(\datapath_1.regfile_1.regOut[2] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

FILL FILL_1__10933_ (
);

BUFX2 BUFX2_insert270 (
    .A(_2379_),
    .Y(_2379__bF$buf2)
);

BUFX2 BUFX2_insert271 (
    .A(_2379_),
    .Y(_2379__bF$buf1)
);

BUFX2 BUFX2_insert272 (
    .A(_2379_),
    .Y(_2379__bF$buf0)
);

BUFX2 BUFX2_insert273 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf4 )
);

BUFX2 BUFX2_insert274 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf3 )
);

AND2X2 _17968_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_6885_)
);

AND2X2 _17548_ (
    .A(_6328__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_6471_)
);

BUFX2 BUFX2_insert275 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf2 )
);

BUFX2 BUFX2_insert276 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf1 )
);

OR2X2 _17128_ (
    .A(_6049_),
    .B(_6056_),
    .Y(_6057_)
);

FILL FILL253840x291460 (
);

BUFX2 BUFX2_insert277 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf0 )
);

BUFX2 BUFX2_insert278 (
    .A(_3605_),
    .Y(_3605__bF$buf4)
);

FILL FILL_0__12398_ (
);

OR2X2 _12683_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(_2247_),
    .Y(_2248_)
);

BUFX2 BUFX2_insert279 (
    .A(_3605_),
    .Y(_3605__bF$buf3)
);

AND2X2 _12263_ (
    .A(_1960_),
    .B(_1959_),
    .Y(_1917_[21])
);

FILL FILL_0__18624_ (
);

FILL FILL50920x227240 (
);

FILL FILL428640x330980 (
);

FILL FILL_0__8725_ (
);

FILL FILL412680x44460 (
);

OR2X2 _13888_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.mux_iord.din0 [24]),
    .Y(_3325_)
);

FILL FILL240160x296400 (
);

AND2X2 _13468_ (
    .A(_3000_),
    .B(_2511_),
    .Y(_3001_)
);

AND2X2 _13048_ (
    .A(_2604_),
    .B(_2310_),
    .Y(_2605_)
);

FILL FILL_1__15971_ (
);

FILL FILL_0__19409_ (
);

FILL FILL_0__14964_ (
);

FILL FILL192280x24700 (
);

FILL FILL_0__14124_ (
);

FILL FILL321480x19760 (
);

FILL FILL_1__11051_ (
);

FILL FILL_0__15749_ (
);

FILL FILL_0__15329_ (
);

AND2X2 _15614_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_4566_)
);

FILL FILL_0__10464_ (
);

AND2X2 _18086_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_7001_)
);

FILL FILL_0__19162_ (
);

FILL FILL88920x167960 (
);

AND2X2 _16819_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_5753_)
);

FILL FILL_0__9683_ (
);

AND2X2 _11954_ (
    .A(_1794_),
    .B(_1793_),
    .Y(_1785_[4])
);

FILL FILL_0__9263_ (
);

DFFSR _11534_ (
    .CLK(clk_bF$buf34),
    .D(_1521_[14]),
    .Q(\datapath_1.regfile_1.regOut[24] [14]),
    .R(rst_bF$buf71),
    .S(vdd)
);

FILL FILL_0__11249_ (
);

AND2X2 _11114_ (
    .A(_1374_),
    .B(_1373_),
    .Y(_1323_[25])
);

FILL FILL128440x256880 (
);

FILL FILL_0__15082_ (
);

INVX1 _12739_ (
    .A(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2304_)
);

DFFSR _12319_ (
    .CLK(clk_bF$buf43),
    .D(_1917_[25]),
    .Q(\datapath_1.regfile_1.regOut[30] [25]),
    .R(rst_bF$buf13),
    .S(vdd)
);

FILL FILL_0__13815_ (
);

FILL FILL_1__17294_ (
);

OR2X2 _16992_ (
    .A(_5922_),
    .B(_5919_),
    .Y(_5923_)
);

AND2X2 _16572_ (
    .A(_4239__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_5509_)
);

OR2X2 _16152_ (
    .A(_5088_),
    .B(_5095_),
    .Y(_5096_)
);

FILL FILL39520x69160 (
);

OR2X2 _8494_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .B(_68__bF$buf4),
    .Y(_28_)
);

FILL FILL_1__10322_ (
);

AND2X2 _17777_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_6697_)
);

AND2X2 _17357_ (
    .A(_6282__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_6283_)
);

FILL FILL_1__19440_ (
);

NOR2X1 _12492_ (
    .A(_2093_),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2095_)
);

OR2X2 _12072_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_1853_)
);

FILL FILL_0__18433_ (
);

FILL FILL_0__18013_ (
);

OR2X2 _9699_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_651_)
);

OR2X2 _9279_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_431_)
);

FILL FILL367840x177840 (
);

FILL FILL_0__8534_ (
);

AND2X2 _10805_ (
    .A(_1208_),
    .B(_1207_),
    .Y(_1191_[8])
);

FILL FILL203680x64220 (
);

AND2X2 _13697_ (
    .A(_3084__bF$buf4),
    .B(\datapath_1.PCJump [15]),
    .Y(_3177_)
);

OR2X2 _13277_ (
    .A(_2219_),
    .B(_2415_),
    .Y(_2820_)
);

FILL FILL67640x187720 (
);

OR2X2 _19503_ (
    .A(gnd),
    .B(_8385__bF$buf1),
    .Y(_8371_)
);

FILL FILL207480x182780 (
);

FILL FILL_0__14773_ (
);

FILL FILL_0__9319_ (
);

FILL FILL335920x311220 (
);

FILL FILL_1__16145_ (
);

FILL FILL_0__15978_ (
);

FILL FILL503120x167960 (
);

OR2X2 _15843_ (
    .A(_4790_),
    .B(_4791_),
    .Y(_4792_)
);

FILL FILL_0__15138_ (
);

AND2X2 _15423_ (
    .A(_4197__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_4378_)
);

DFFSR _15003_ (
    .CLK(clk_bF$buf12),
    .D(_3936_[22]),
    .Q(\datapath_1.mux_iord.din0 [22]),
    .R(rst_bF$buf5),
    .S(vdd)
);

FILL FILL_0__10693_ (
);

FILL FILL_0__10273_ (
);

FILL FILL344280x108680 (
);

FILL FILL147440x370500 (
);

FILL FILL_0__19391_ (
);

AND2X2 _16628_ (
    .A(_4225__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_5565_)
);

OR2X2 _16208_ (
    .A(_5147_),
    .B(_5150_),
    .Y(_5151_)
);

FILL FILL_0__9492_ (
);

FILL FILL_0__11898_ (
);

OR2X2 _11763_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_1707_)
);

FILL FILL_0__11058_ (
);

OR2X2 _11343_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_1487_)
);

FILL FILL_0__17704_ (
);

FILL FILL164160x286520 (
);

FILL FILL121600x182780 (
);

AND2X2 _9911_ (
    .A(_752_),
    .B(_751_),
    .Y(_729_[11])
);

OR2X2 _12968_ (
    .A(_2157__bF$buf2),
    .B(_2529_),
    .Y(_2530_)
);

FILL FILL_1_BUFX2_insert982 (
);

OR2X2 _12548_ (
    .A(_2125_),
    .B(_2136_),
    .Y(_2137_)
);

AND2X2 _12128_ (
    .A(_1890_),
    .B(_1889_),
    .Y(_1851_[19])
);

FILL FILL_1_BUFX2_insert984 (
);

FILL FILL_1_BUFX2_insert986 (
);

FILL FILL_0__18909_ (
);

FILL FILL_0__13624_ (
);

FILL FILL65360x370500 (
);

FILL FILL356440x335920 (
);

FILL FILL_0__16096_ (
);

OR2X2 _16381_ (
    .A(_5319_),
    .B(_5320_),
    .Y(_5321_)
);

FILL FILL300200x370500 (
);

FILL FILL_1__9653_ (
);

FILL FILL310080x316160 (
);

FILL FILL373920x345800 (
);

FILL FILL_0__14829_ (
);

FILL FILL_0__14409_ (
);

BUFX2 BUFX2_insert650 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf4 )
);

BUFX2 BUFX2_insert651 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf3 )
);

BUFX2 BUFX2_insert652 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf2 )
);

FILL FILL375440x44460 (
);

BUFX2 BUFX2_insert653 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf1 )
);

FILL FILL82080x286520 (
);

BUFX2 BUFX2_insert654 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf0 )
);

OR2X2 _17586_ (
    .A(_6500_),
    .B(_6508_),
    .Y(_6509_)
);

BUFX2 BUFX2_insert655 (
    .A(_4154_),
    .Y(_4154__bF$buf4)
);

BUFX2 BUFX2_insert656 (
    .A(_4154_),
    .Y(_4154__bF$buf3)
);

AND2X2 _17166_ (
    .A(_4167__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_6094_)
);

BUFX2 BUFX2_insert657 (
    .A(_4154_),
    .Y(_4154__bF$buf2)
);

BUFX2 BUFX2_insert658 (
    .A(_4154_),
    .Y(_4154__bF$buf1)
);

BUFX2 BUFX2_insert659 (
    .A(_4154_),
    .Y(_4154__bF$buf0)
);

FILL FILL_0__18662_ (
);

FILL FILL_0__18242_ (
);

FILL FILL76000x242060 (
);

FILL FILL409640x237120 (
);

DFFSR _9088_ (
    .CLK(clk_bF$buf19),
    .D(_267_[19]),
    .Q(\datapath_1.regfile_1.regOut[5] [19]),
    .R(rst_bF$buf13),
    .S(vdd)
);

FILL FILL_0__8763_ (
);

FILL FILL53960x143260 (
);

OR2X2 _10614_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_1121_)
);

FILL FILL445360x9880 (
);

FILL FILL285000x113620 (
);

NAND2X1 _13086_ (
    .A(_2467_),
    .B(_2379__bF$buf0),
    .Y(_2641_)
);

FILL FILL_0__19027_ (
);

AND2X2 _19312_ (
    .A(_6244__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_8208_)
);

FILL FILL_0__14582_ (
);

FILL FILL431680x340860 (
);

FILL FILL266000x271700 (
);

FILL FILL_0__9968_ (
);

FILL FILL_0__9548_ (
);

FILL FILL_0__9128_ (
);

AND2X2 _11819_ (
    .A(_1724_),
    .B(_1723_),
    .Y(_1719_[2])
);

FILL FILL348840x350740 (
);

FILL FILL_1__16794_ (
);

FILL FILL_1__16374_ (
);

FILL FILL_0__15367_ (
);

AND2X2 _15652_ (
    .A(_4236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_4604_)
);

AND2X2 _15232_ (
    .A(_4189__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_4190_)
);

FILL FILL_0__10082_ (
);

FILL FILL_1__8924_ (
);

FILL FILL114760x163020 (
);

FILL FILL_1__17159_ (
);

OR2X2 _16857_ (
    .A(_5774_),
    .B(_5789_),
    .Y(_5790_)
);

OR2X2 _16437_ (
    .A(_5376_),
    .B(_5375_),
    .Y(_5377_)
);

AND2X2 _16017_ (
    .A(_4217__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_4963_)
);

OR2X2 _11992_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .B(_1850__bF$buf0),
    .Y(_1820_)
);

OR2X2 _11572_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .B(_1652__bF$buf1),
    .Y(_1600_)
);

DFFSR _11152_ (
    .CLK(clk_bF$buf81),
    .D(_1323_[19]),
    .Q(\datapath_1.regfile_1.regOut[21] [19]),
    .R(rst_bF$buf19),
    .S(vdd)
);

FILL FILL498560x222300 (
);

FILL FILL_0__17933_ (
);

FILL FILL_0__17513_ (
);

OR2X2 _8779_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .B(_200__bF$buf4),
    .Y(_178_)
);

DFFSR _9720_ (
    .CLK(clk_bF$buf59),
    .D(_597_[6]),
    .Q(\datapath_1.regfile_1.regOut[10] [6]),
    .R(rst_bF$buf92),
    .S(vdd)
);

OR2X2 _9300_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_445_)
);

FILL FILL_1__13499_ (
);

FILL FILL337440x74100 (
);

AND2X2 _12777_ (
    .A(_2339_),
    .B(_2341_),
    .Y(_2342_)
);

FILL FILL_1__19305_ (
);

OR2X2 _12357_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_2003_)
);

FILL FILL269800x49400 (
);

FILL FILL_1__14440_ (
);

FILL FILL_0__13433_ (
);

FILL FILL_0__13013_ (
);

FILL FILL131480x266760 (
);

AND2X2 _16190_ (
    .A(_4203__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_5133_)
);

FILL FILL_1__9042_ (
);

FILL FILL_1__10780_ (
);

FILL FILL_0__14638_ (
);

AND2X2 _14923_ (
    .A(_3961_),
    .B(_3960_),
    .Y(_3936_[12])
);

FILL FILL_0__14218_ (
);

AND2X2 _14503_ (
    .A(_3741_),
    .B(_3740_),
    .Y(_3738_[1])
);

FILL FILL355680x103740 (
);

FILL FILL183160x14820 (
);

AND2X2 _17395_ (
    .A(_6258_),
    .B(_6209_),
    .Y(_6321_)
);

FILL FILL_0__18891_ (
);

FILL FILL152760x197600 (
);

FILL FILL_1__11985_ (
);

OR2X2 _15708_ (
    .A(_4658_),
    .B(_4657_),
    .Y(_4659_)
);

FILL FILL_0__10978_ (
);

OR2X2 _10843_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_1256__bF$buf1),
    .Y(_1234_)
);

OR2X2 _10423_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .B(_1058__bF$buf4),
    .Y(_1014_)
);

DFFSR _10003_ (
    .CLK(clk_bF$buf10),
    .D(_729_[31]),
    .Q(\datapath_1.regfile_1.regOut[12] [31]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _19541_ (
    .CLK(clk_bF$buf63),
    .D(_8320_[18]),
    .Q(\datapath_1.regfile_1.regOut[0] [18]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL_0__19256_ (
);

AND2X2 _19121_ (
    .A(_6236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_8020_)
);

FILL FILL_0__14391_ (
);

FILL FILL152000x321100 (
);

FILL FILL_0__9777_ (
);

OR2X2 _11628_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_1637_)
);

OR2X2 _11208_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_1417_)
);

FILL FILL_1__13711_ (
);

FILL FILL_0__15596_ (
);

OR2X2 _15881_ (
    .A(_4828_),
    .B(_4821_),
    .Y(_4829_)
);

AND2X2 _15461_ (
    .A(_4225__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_4416_)
);

INVX1 _15041_ (
    .A(_4006_),
    .Y(_4030_)
);

FILL FILL_1__8733_ (
);

FILL FILL416480x217360 (
);

FILL FILL449920x9880 (
);

FILL FILL_0__13909_ (
);

FILL FILL19000x276640 (
);

AND2X2 _16666_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_5602_)
);

FILL FILL237120x172900 (
);

OR2X2 _16246_ (
    .A(_5185_),
    .B(_5188_),
    .Y(_5189_)
);

AND2X2 _11381_ (
    .A(_1512_),
    .B(_1511_),
    .Y(_1455_[28])
);

FILL FILL_0__11096_ (
);

FILL FILL_1__9938_ (
);

FILL FILL186200x340860 (
);

FILL FILL433960x227240 (
);

FILL FILL439280x301340 (
);

FILL FILL_0__17742_ (
);

AND2X2 _8588_ (
    .A(_70_),
    .B(_133_),
    .Y(_69_[0])
);

FILL FILL219640x345800 (
);

DFFSR _12586_ (
    .CLK(clk_bF$buf23),
    .D(_2143_[2]),
    .Q(\control_1.reg_state.dout [2]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _12166_ (
    .CLK(clk_bF$buf4),
    .D(_1851_[1]),
    .Q(\datapath_1.regfile_1.regOut[29] [1]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _18812_ (
    .A(_7715_),
    .B(_7714_),
    .Y(_7716_)
);

FILL FILL_0__18527_ (
);

FILL FILL_0__18107_ (
);

FILL FILL_0__13662_ (
);

FILL FILL_0__13242_ (
);

FILL FILL_0__8628_ (
);

FILL FILL268280x370500 (
);

FILL FILL126920x29640 (
);

DFFSR _14732_ (
    .CLK(clk_bF$buf80),
    .D(_3804_[9]),
    .Q(\datapath_1.a [9]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__14447_ (
);

OR2X2 _14312_ (
    .A(vdd),
    .B(ALUOut[24]),
    .Y(_3654_)
);

CLKBUF1 CLKBUF1_insert190 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert191 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert192 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert193 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert194 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert195 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert196 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert197 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert198 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert199 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf24)
);

FILL FILL148200x123500 (
);

FILL FILL_0__18280_ (
);

FILL FILL30400x227240 (
);

FILL FILL_1__16659_ (
);

FILL FILL_1__16239_ (
);

FILL FILL_1__11374_ (
);

OR2X2 _15937_ (
    .A(_4883_),
    .B(_4880_),
    .Y(_4884_)
);

AND2X2 _15517_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_4471_)
);

FILL FILL_0__10787_ (
);

FILL FILL_1__17600_ (
);

AND2X2 _10652_ (
    .A(_1126_),
    .B(_1189_),
    .Y(_1125_[0])
);

DFFSR _10232_ (
    .CLK(clk_bF$buf51),
    .D(_861_[2]),
    .Q(\datapath_1.regfile_1.regOut[14] [2]),
    .R(rst_bF$buf52),
    .S(vdd)
);

FILL FILL_0__19485_ (
);

FILL FILL_0__19065_ (
);

AND2X2 _19350_ (
    .A(_6315__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_8246_)
);

OR2X2 _8800_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .B(_200__bF$buf1),
    .Y(_192_)
);

FILL FILL_1__12999_ (
);

FILL FILL_0__9166_ (
);

OR2X2 _11857_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .B(_1784__bF$buf4),
    .Y(_1750_)
);

OR2X2 _11437_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .B(_1586__bF$buf2),
    .Y(_1530_)
);

DFFSR _11017_ (
    .CLK(clk_bF$buf47),
    .D(_1257_[13]),
    .Q(\datapath_1.regfile_1.regOut[20] [13]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL_1__13940_ (
);

FILL FILL348080x326040 (
);

FILL FILL228760x276640 (
);

FILL FILL_0__12933_ (
);

FILL FILL_0__12513_ (
);

FILL FILL192280x316160 (
);

AND2X2 _15690_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_4641_)
);

AND2X2 _15270_ (
    .A(_4222_),
    .B(_4144_),
    .Y(_4228_)
);

FILL FILL409640x54340 (
);

FILL FILL161880x29640 (
);

FILL FILL_0__13718_ (
);

FILL FILL22800x242060 (
);

FILL FILL117800x83980 (
);

AND2X2 _16895_ (
    .A(_4177__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_5827_)
);

AND2X2 _16475_ (
    .A(_4151__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_5414_)
);

OR2X2 _16055_ (
    .A(_4993_),
    .B(_5000_),
    .Y(_5001_)
);

OR2X2 _11190_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_1405_)
);

FILL FILL_1__9747_ (
);

FILL FILL_0__17551_ (
);

FILL FILL_0__17131_ (
);

FILL FILL22040x29640 (
);

BUFX2 _8397_ (
    .A(_1_[5]),
    .Y(memoryAddress[5])
);

FILL FILL469680x350740 (
);

FILL FILL125400x266760 (
);

AND2X2 _12395_ (
    .A(_2028_),
    .B(_2027_),
    .Y(_1983_[22])
);

FILL FILL_0__18756_ (
);

OR2X2 _18621_ (
    .A(_7526_),
    .B(_7527_),
    .Y(_7528_)
);

FILL FILL294880x177840 (
);

AND2X2 _18201_ (
    .A(_6289__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_7114_)
);

FILL FILL_0__13891_ (
);

FILL FILL_0__13471_ (
);

FILL FILL_0__8857_ (
);

OR2X2 _10708_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .B(_1190__bF$buf3),
    .Y(_1164_)
);

FILL FILL_1__15263_ (
);

OR2X2 _19406_ (
    .A(_8293_),
    .B(_8300_),
    .Y(_8301_)
);

OR2X2 _14961_ (
    .A(\datapath_1.mux_pcsrc.dout [25]),
    .B(_4001__bF$buf2),
    .Y(_3987_)
);

FILL FILL_0__14256_ (
);

OR2X2 _14541_ (
    .A(memoryOutData[14]),
    .B(_3803__bF$buf2),
    .Y(_3767_)
);

AND2X2 _14121_ (
    .A(_3344__bF$buf1),
    .B(gnd),
    .Y(_3523_)
);

FILL FILL207480x296400 (
);

FILL FILL53960x306280 (
);

FILL FILL357960x217360 (
);

FILL FILL_1__16888_ (
);

FILL FILL6080x9880 (
);

FILL FILL_1__11183_ (
);

AND2X2 _15746_ (
    .A(_4158__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_4696_)
);

AND2X2 _15326_ (
    .A(_4172__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_4283_)
);

FILL FILL_0__10596_ (
);

DFFSR _10881_ (
    .CLK(clk_bF$buf49),
    .D(_1191_[6]),
    .Q(\datapath_1.regfile_1.regOut[19] [6]),
    .R(rst_bF$buf66),
    .S(vdd)
);

OR2X2 _10461_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_1039_)
);

OR2X2 _10041_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_819_)
);

FILL FILL_0__16822_ (
);

FILL FILL_0__16402_ (
);

FILL FILL275880x123500 (
);

FILL FILL243960x335920 (
);

FILL FILL_0__9395_ (
);

DFFSR _11666_ (
    .CLK(clk_bF$buf8),
    .D(_1587_[17]),
    .Q(\datapath_1.regfile_1.regOut[25] [17]),
    .R(rst_bF$buf10),
    .S(vdd)
);

AND2X2 _11246_ (
    .A(_1442_),
    .B(_1441_),
    .Y(_1389_[26])
);

FILL FILL_0__17607_ (
);

FILL FILL186960x286520 (
);

FILL FILL_0__12742_ (
);

OR2X2 _9814_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .B(_728__bF$buf4),
    .Y(_708_)
);

FILL FILL_1__14114_ (
);

FILL FILL_0__13947_ (
);

AND2X2 _13812_ (
    .A(_3089__bF$buf1),
    .B(gnd),
    .Y(_3276_)
);

FILL FILL_0__13107_ (
);

FILL FILL422560x182780 (
);

FILL FILL319960x321100 (
);

OR2X2 _16284_ (
    .A(_5224_),
    .B(_5225_),
    .Y(_5226_)
);

FILL FILL332880x316160 (
);

FILL FILL_0__17780_ (
);

FILL FILL_0__17360_ (
);

FILL FILL_1__15739_ (
);

FILL FILL_1__10874_ (
);

FILL FILL22040x286520 (
);

OR2X2 _17489_ (
    .A(_6412_),
    .B(_6411_),
    .Y(_6413_)
);

AND2X2 _17069_ (
    .A(_4223__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_5999_)
);

FILL FILL273600x29640 (
);

OR2X2 _18850_ (
    .A(_7752_),
    .B(_7751_),
    .Y(_7753_)
);

FILL FILL_0__18145_ (
);

OR2X2 _18430_ (
    .A(_7339_),
    .B(_7335_),
    .Y(_7340_)
);

FILL FILL180880x227240 (
);

OR2X2 _18010_ (
    .A(_6925_),
    .B(_6918_),
    .Y(_6926_)
);

FILL FILL88160x29640 (
);

FILL FILL170240x187720 (
);

FILL FILL_0__8666_ (
);

AND2X2 _10937_ (
    .A(_1276_),
    .B(_1275_),
    .Y(_1257_[9])
);

DFFSR _10517_ (
    .CLK(clk_bF$buf8),
    .D(_993_[29]),
    .Q(\datapath_1.regfile_1.regOut[16] [29]),
    .R(rst_bF$buf77),
    .S(vdd)
);

FILL FILL_1__15492_ (
);

FILL FILL129200x306280 (
);

AND2X2 _19215_ (
    .A(_6289__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_8113_)
);

AND2X2 _14770_ (
    .A(_3879_),
    .B(_3878_),
    .Y(_3870_[4])
);

FILL FILL_0__14065_ (
);

DFFSR _14350_ (
    .CLK(clk_bF$buf62),
    .D(_3606_[14]),
    .Q(ALUOut[14]),
    .R(rst_bF$buf18),
    .S(vdd)
);

FILL FILL275880x24700 (
);

FILL FILL_1__13805_ (
);

OR2X2 _15975_ (
    .A(_4918_),
    .B(_4921_),
    .Y(_4922_)
);

AND2X2 _15555_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_4508_)
);

NOR2X1 _15135_ (
    .A(_4060_),
    .B(_4042_),
    .Y(\datapath_1.regfile_1.regEn [18])
);

OR2X2 _10690_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_1190__bF$buf3),
    .Y(_1152_)
);

OR2X2 _10270_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .B(_992__bF$buf4),
    .Y(_932_)
);

FILL FILL_0__16631_ (
);

FILL FILL_0__16211_ (
);

OR2X2 _11895_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .Y(_1775_)
);

FILL FILL_1__18423_ (
);

OR2X2 _11475_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_1555_)
);

OR2X2 _11055_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_1335_)
);

FILL FILL_1__18003_ (
);

AND2X2 _17701_ (
    .A(_6282__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_6622_)
);

FILL FILL279680x24700 (
);

FILL FILL_0__12131_ (
);

FILL FILL449920x291460 (
);

AND2X2 _9623_ (
    .A(_600_),
    .B(_599_),
    .Y(_597_[1])
);

DFFSR _9203_ (
    .CLK(clk_bF$buf70),
    .D(_333_[5]),
    .Q(\datapath_1.regfile_1.regOut[6] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

FILL FILL269040x123500 (
);

FILL FILL28880x128440 (
);

AND2X2 _18906_ (
    .A(_6206__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_7808_)
);

FILL FILL208240x232180 (
);

FILL FILL_0__13756_ (
);

FILL FILL_0__13336_ (
);

OR2X2 _13621_ (
    .A(_3110_),
    .B(_3111_),
    .Y(_3112_)
);

OR2X2 _13201_ (
    .A(_2387__bF$buf3),
    .B(_2749_),
    .Y(_2750_)
);

AND2X2 _16093_ (
    .A(_4236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_5038_)
);

FILL FILL472720x148200 (
);

FILL FILL_1__9785_ (
);

FILL FILL_1__15128_ (
);

FILL FILL_1__10683_ (
);

OR2X2 _14826_ (
    .A(\datapath_1.rd2 [23]),
    .B(_3935__bF$buf4),
    .Y(_3917_)
);

OR2X2 _14406_ (
    .A(memoryOutData[12]),
    .B(_3737__bF$buf1),
    .Y(_3697_)
);

OR2X2 _17298_ (
    .A(_6213_),
    .B(_6223_),
    .Y(_6224_)
);

FILL FILL470440x93860 (
);

FILL FILL132240x74100 (
);

FILL FILL_0__15902_ (
);

FILL FILL_0__18794_ (
);

FILL FILL_0__18374_ (
);

FILL FILL294120x345800 (
);

FILL FILL_0__8475_ (
);

DFFSR _10746_ (
    .CLK(clk_bF$buf19),
    .D(_1125_[0]),
    .Q(\datapath_1.regfile_1.regOut[18] [0]),
    .R(rst_bF$buf79),
    .S(vdd)
);

OR2X2 _10326_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_969_)
);

FILL FILL12920x123500 (
);

FILL FILL_0__11822_ (
);

FILL FILL229520x350740 (
);

AND2X2 _19444_ (
    .A(_8331_),
    .B(_8330_),
    .Y(_8320_[5])
);

AND2X2 _19024_ (
    .A(_6250__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_7925_)
);

FILL FILL_0__12607_ (
);

FILL FILL_1_BUFX2_insert225 (
);

FILL FILL_1_BUFX2_insert227 (
);

FILL FILL246240x266760 (
);

OR2X2 _15784_ (
    .A(_4726_),
    .B(_4733_),
    .Y(_4734_)
);

FILL FILL_0__15499_ (
);

OR2X2 _15364_ (
    .A(_4319_),
    .B(_4318_),
    .Y(_4320_)
);

FILL FILL_0__15079_ (
);

FILL FILL_1__8636_ (
);

FILL FILL_0__16860_ (
);

FILL FILL_0__16020_ (
);

FILL FILL_1__14819_ (
);

AND2X2 _16989_ (
    .A(_4175__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_5920_)
);

OR2X2 _16569_ (
    .A(_5475_),
    .B(_5506_),
    .Y(_5507_)
);

AND2X2 _16149_ (
    .A(_4151__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_5093_)
);

FILL FILL_1__18652_ (
);

DFFSR _11284_ (
    .CLK(clk_bF$buf25),
    .D(_1389_[22]),
    .Q(\datapath_1.regfile_1.regOut[22] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

FILL FILL487920x113620 (
);

FILL FILL112480x69160 (
);

AND2X2 _17930_ (
    .A(_6847_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.rd1 [8])
);

FILL FILL_0__17645_ (
);

FILL FILL464360x256880 (
);

FILL FILL_0__17225_ (
);

AND2X2 _17510_ (
    .A(_6255__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_6434_)
);

FILL FILL_0__12780_ (
);

DFFSR _9852_ (
    .CLK(clk_bF$buf75),
    .D(_663_[9]),
    .Q(\datapath_1.regfile_1.regOut[11] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

OR2X2 _9432_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_513_)
);

OR2X2 _9012_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_293_)
);

NAND3X1 _12489_ (
    .A(_2092_),
    .B(\control_1.reg_state.dout [3]),
    .C(_2093_),
    .Y(_2094_)
);

FILL FILL310080x202540 (
);

INVX2 _12069_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .Y(_1916_)
);

FILL FILL_1__14152_ (
);

NOR2X1 _18715_ (
    .A(_6310__bF$buf3),
    .B(_7619_),
    .Y(_7620_)
);

FILL FILL_0__13985_ (
);

OR2X2 _13850_ (
    .A(\datapath_1.a [11]),
    .B(_3342__bF$buf3),
    .Y(_3300_)
);

XNOR2X1 _13430_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2964_)
);

AND2X2 _13010_ (
    .A(_2569_),
    .B(_2567_),
    .Y(_2570_)
);

FILL FILL194560x74100 (
);

FILL FILL253080x153140 (
);

FILL FILL323760x69160 (
);

FILL FILL_1__15777_ (
);

FILL FILL_1__15357_ (
);

FILL FILL_1__10072_ (
);

AND2X2 _14635_ (
    .A(_3809_),
    .B(_3808_),
    .Y(_3804_[2])
);

OR2X2 _14215_ (
    .A(MemToReg_bF$buf4),
    .B(ALUOut[24]),
    .Y(_3588_)
);

FILL FILL445360x202540 (
);

FILL FILL_0__18183_ (
);

FILL FILL242440x296400 (
);

OR2X2 _10975_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .B(_1322__bF$buf1),
    .Y(_1302_)
);

OR2X2 _10555_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .B(_1124__bF$buf2),
    .Y(_1082_)
);

OR2X2 _10135_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(_926__bF$buf0),
    .Y(_862_)
);

FILL FILL_0__16916_ (
);

FILL FILL449160x123500 (
);

FILL FILL_0__11211_ (
);

NOR2X1 _19253_ (
    .A(_6310__bF$buf2),
    .B(_8149_),
    .Y(_8150_)
);

DFFSR _8703_ (
    .CLK(clk_bF$buf43),
    .D(_69_[21]),
    .Q(\datapath_1.regfile_1.regOut[2] [21]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL56240x375440 (
);

FILL FILL_0__9489_ (
);

FILL FILL_0__12836_ (
);

OR2X2 _12701_ (
    .A(\datapath_1.alu_1.ALUInA [23]),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2266_)
);

FILL FILL_0__12416_ (
);

FILL FILL119320x321100 (
);

AND2X2 _15593_ (
    .A(_4234__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_4546_)
);

AND2X2 _15173_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_4131_)
);

AND2X2 _9908_ (
    .A(_750_),
    .B(_749_),
    .Y(_729_[10])
);

FILL FILL_1__8445_ (
);

FILL FILL200640x54340 (
);

FILL FILL_1__14628_ (
);

OR2X2 _13906_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.PCJump [30]),
    .Y(_3337_)
);

AND2X2 _16798_ (
    .A(_4175__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_5732_)
);

AND2X2 _16378_ (
    .A(_5318_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd2 [17])
);

AND2X2 _11093_ (
    .A(_1360_),
    .B(_1359_),
    .Y(_1323_[18])
);

FILL FILL_1__18041_ (
);

FILL FILL_0__17874_ (
);

FILL FILL236360x330980 (
);

FILL FILL_1__10968_ (
);

OR2X2 _9661_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .B(_662__bF$buf3),
    .Y(_626_)
);

OR2X2 _9241_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_464__bF$buf3),
    .Y(_406_)
);

DFFSR _12298_ (
    .CLK(clk_bF$buf87),
    .D(_1917_[4]),
    .Q(\datapath_1.regfile_1.regOut[30] [4]),
    .R(rst_bF$buf2),
    .S(vdd)
);

FILL FILL_0__18659_ (
);

AND2X2 _18944_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_7846_)
);

FILL FILL_0__18239_ (
);

AND2X2 _18524_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_7432_)
);

OR2X2 _18104_ (
    .A(_7018_),
    .B(_7017_),
    .Y(_7019_)
);

FILL FILL_0__13374_ (
);

FILL FILL196840x291460 (
);

OR2X2 _19309_ (
    .A(_8203_),
    .B(_8204_),
    .Y(_8205_)
);

FILL FILL71440x247000 (
);

DFFSR _14864_ (
    .CLK(clk_bF$buf58),
    .D(_3870_[12]),
    .Q(_2_[12]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__14159_ (
);

OR2X2 _14444_ (
    .A(vdd),
    .B(\datapath_1.Data [25]),
    .Y(_3722_)
);

AND2X2 _14024_ (
    .A(_3347__bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3440_)
);

FILL FILL161120x34580 (
);

FILL FILL_0__15940_ (
);

FILL FILL452960x167960 (
);

FILL FILL_0__15520_ (
);

FILL FILL_0__15100_ (
);

FILL FILL226480x64220 (
);

AND2X2 _15649_ (
    .A(_4158__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [6]),
    .Y(_4601_)
);

AND2X2 _15229_ (
    .A(_4186_),
    .B(_4144_),
    .Y(_4187_)
);

AND2X2 _10784_ (
    .A(_1194_),
    .B(_1193_),
    .Y(_1191_[1])
);

FILL FILL_0__10079_ (
);

DFFSR _10364_ (
    .CLK(clk_bF$buf66),
    .D(_927_[5]),
    .Q(\datapath_1.regfile_1.regOut[15] [5]),
    .R(rst_bF$buf80),
    .S(vdd)
);

FILL FILL69920x187720 (
);

FILL FILL_0__16725_ (
);

FILL FILL209760x182780 (
);

FILL FILL_0__11860_ (
);

FILL FILL_0__19197_ (
);

OR2X2 _19482_ (
    .A(gnd),
    .B(_8385__bF$buf2),
    .Y(_8357_)
);

OR2X2 _19062_ (
    .A(_7961_),
    .B(_7960_),
    .Y(_7962_)
);

OR2X2 _8932_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .B(_266__bF$buf1),
    .Y(_260_)
);

OR2X2 _8512_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .B(_68__bF$buf1),
    .Y(_40_)
);

FILL FILL_0__9298_ (
);

FILL FILL_1__18937_ (
);

OR2X2 _11989_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_1850__bF$buf0),
    .Y(_1818_)
);

FILL FILL_1__18517_ (
);

OR2X2 _11569_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .B(_1652__bF$buf1),
    .Y(_1598_)
);

DFFSR _11149_ (
    .CLK(clk_bF$buf64),
    .D(_1323_[16]),
    .Q(\datapath_1.regfile_1.regOut[21] [16]),
    .R(rst_bF$buf10),
    .S(vdd)
);

FILL FILL_1__13232_ (
);

FILL FILL269040x4940 (
);

FILL FILL505400x167960 (
);

AND2X2 _12930_ (
    .A(_2494_),
    .B(_2373_),
    .Y(_2495_)
);

FILL FILL_0__12225_ (
);

NAND2X1 _12510_ (
    .A(\control_1.reg_state.dout [3]),
    .B(_2093_),
    .Y(_2105_)
);

FILL FILL_1_BUFX2_insert603 (
);

FILL FILL_1_BUFX2_insert605 (
);

FILL FILL_1_BUFX2_insert607 (
);

FILL FILL346560x108680 (
);

FILL FILL97280x69160 (
);

DFFSR _9717_ (
    .CLK(clk_bF$buf56),
    .D(_597_[3]),
    .Q(\datapath_1.regfile_1.regOut[10] [3]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL457520x79040 (
);

FILL FILL288040x4940 (
);

OR2X2 _13715_ (
    .A(_3192_),
    .B(_3191_),
    .Y(_3193_)
);

AND2X2 _16187_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_5130_)
);

FILL FILL_1__9879_ (
);

FILL FILL_0__17263_ (
);

FILL FILL330600x64220 (
);

AND2X2 _9890_ (
    .A(_738_),
    .B(_737_),
    .Y(_729_[4])
);

DFFSR _9470_ (
    .CLK(clk_bF$buf63),
    .D(_465_[14]),
    .Q(\datapath_1.regfile_1.regOut[8] [14]),
    .R(rst_bF$buf7),
    .S(vdd)
);

AND2X2 _9050_ (
    .A(_318_),
    .B(_317_),
    .Y(_267_[25])
);

FILL FILL77520x39520 (
);

FILL FILL367080x266760 (
);

FILL FILL505400x74100 (
);

FILL FILL_0__18888_ (
);

FILL FILL358720x335920 (
);

AND2X2 _18753_ (
    .A(_6264__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_7658_)
);

FILL FILL_0__18468_ (
);

AND2X2 _18333_ (
    .A(_6302__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_7244_)
);

FILL FILL_0__18048_ (
);

FILL FILL80560x365560 (
);

FILL FILL_0__13183_ (
);

FILL FILL_0__8989_ (
);

FILL FILL312360x316160 (
);

FILL FILL_1__12923_ (
);

FILL FILL_1__12503_ (
);

FILL FILL_0__9930_ (
);

FILL FILL398240x44460 (
);

DFFSR _19538_ (
    .CLK(clk_bF$buf104),
    .D(_8320_[15]),
    .Q(\datapath_1.regfile_1.regOut[0] [15]),
    .R(rst_bF$buf80),
    .S(vdd)
);

FILL FILL84360x286520 (
);

AND2X2 _19118_ (
    .A(_6250__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_8017_)
);

OR2X2 _14673_ (
    .A(\datapath_1.rd1 [15]),
    .B(_3869__bF$buf0),
    .Y(_3835_)
);

OR2X2 _14253_ (
    .A(\datapath_1.ALUResult [4]),
    .B(_3671__bF$buf2),
    .Y(_3615_)
);

FILL FILL64600x93860 (
);

AND2X2 _15878_ (
    .A(_4183__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_4826_)
);

AND2X2 _15458_ (
    .A(_4236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_4413_)
);

AND2X2 _15038_ (
    .A(_4021_),
    .B(_4026_),
    .Y(_4027_)
);

FILL FILL_1__17541_ (
);

OR2X2 _10593_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_1107_)
);

OR2X2 _10173_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_887_)
);

FILL FILL_1__17121_ (
);

FILL FILL278920x311220 (
);

FILL FILL348080x212420 (
);

FILL FILL437000x276640 (
);

FILL FILL_0__16114_ (
);

FILL FILL433960x340860 (
);

OR2X2 _19291_ (
    .A(_8180_),
    .B(_8187_),
    .Y(_8188_)
);

AND2X2 _8741_ (
    .A(_152_),
    .B(_151_),
    .Y(_135_[8])
);

DFFSR _11798_ (
    .CLK(clk_bF$buf46),
    .D(_1653_[20]),
    .Q(\datapath_1.regfile_1.regOut[26] [20]),
    .R(rst_bF$buf97),
    .S(vdd)
);

AND2X2 _11378_ (
    .A(_1510_),
    .B(_1509_),
    .Y(_1455_[27])
);

FILL FILL_1__13881_ (
);

FILL FILL376960x291460 (
);

FILL FILL_0__17739_ (
);

OR2X2 _17604_ (
    .A(_6492_),
    .B(_6526_),
    .Y(_6527_)
);

FILL FILL_0__17319_ (
);

FILL FILL503120x98800 (
);

FILL FILL_0__12874_ (
);

FILL FILL_0__12034_ (
);

OR2X2 _9946_ (
    .A(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .B(_794__bF$buf1),
    .Y(_776_)
);

OR2X2 _9526_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .B(_596__bF$buf0),
    .Y(_556_)
);

OR2X2 _9106_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .B(_398__bF$buf4),
    .Y(_336_)
);

FILL FILL_1__8483_ (
);

FILL FILL181640x345800 (
);

FILL FILL_1__14246_ (
);

OR2X2 _18809_ (
    .A(_7711_),
    .B(_7712_),
    .Y(_7713_)
);

FILL FILL_0_BUFX2_insert260 (
);

FILL FILL363280x296400 (
);

FILL FILL13680x232180 (
);

FILL FILL_0_BUFX2_insert262 (
);

OR2X2 _13944_ (
    .A(_3371_),
    .B(_3370_),
    .Y(_3372_)
);

FILL FILL_0_BUFX2_insert264 (
);

FILL FILL_0__13239_ (
);

AND2X2 _13524_ (
    .A(_3037_),
    .B(_3036_),
    .Y(_1_[11])
);

NAND2X1 _13104_ (
    .A(_2274_),
    .B(_2504_),
    .Y(_2658_)
);

FILL FILL_0_BUFX2_insert266 (
);

FILL FILL_0_BUFX2_insert267 (
);

FILL FILL_0_BUFX2_insert268 (
);

FILL FILL_0_BUFX2_insert269 (
);

FILL FILL95760x330980 (
);

FILL FILL_1__9688_ (
);

FILL FILL418000x222300 (
);

BUFX2 BUFX2_insert1180 (
    .A(rst),
    .Y(rst_hier0_bF$buf9)
);

BUFX2 BUFX2_insert1181 (
    .A(rst),
    .Y(rst_hier0_bF$buf8)
);

FILL FILL_0__17492_ (
);

BUFX2 BUFX2_insert1182 (
    .A(rst),
    .Y(rst_hier0_bF$buf7)
);

FILL FILL_0__17072_ (
);

BUFX2 BUFX2_insert1183 (
    .A(rst),
    .Y(rst_hier0_bF$buf6)
);

BUFX2 BUFX2_insert1184 (
    .A(rst),
    .Y(rst_hier0_bF$buf5)
);

FILL FILL222680x103740 (
);

BUFX2 BUFX2_insert1185 (
    .A(rst),
    .Y(rst_hier0_bF$buf4)
);

BUFX2 BUFX2_insert1186 (
    .A(rst),
    .Y(rst_hier0_bF$buf3)
);

BUFX2 BUFX2_insert1187 (
    .A(rst),
    .Y(rst_hier0_bF$buf2)
);

BUFX2 BUFX2_insert1188 (
    .A(rst),
    .Y(rst_hier0_bF$buf1)
);

BUFX2 BUFX2_insert1189 (
    .A(rst),
    .Y(rst_hier0_bF$buf0)
);

DFFSR _14729_ (
    .CLK(clk_bF$buf80),
    .D(_3804_[6]),
    .Q(\datapath_1.a [6]),
    .R(rst_bF$buf104),
    .S(vdd)
);

OR2X2 _14309_ (
    .A(vdd),
    .B(ALUOut[23]),
    .Y(_3652_)
);

FILL FILL_0__15805_ (
);

FILL FILL_0__10940_ (
);

FILL FILL_0__10520_ (
);

FILL FILL_0__10100_ (
);

FILL FILL370880x232180 (
);

FILL FILL_0__18697_ (
);

AND2X2 _18982_ (
    .A(_6238__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_7883_)
);

AND2X2 _18562_ (
    .A(_6293__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_7470_)
);

AND2X2 _18142_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_7056_)
);

FILL FILL139080x340860 (
);

FILL FILL270560x326040 (
);

FILL FILL_0__8798_ (
);

OR2X2 _10649_ (
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .Y(_1189_)
);

AND2X2 _10229_ (
    .A(_924_),
    .B(_923_),
    .Y(_861_[31])
);

FILL FILL357960x103740 (
);

FILL FILL_0__11725_ (
);

FILL FILL_0__11305_ (
);

OR2X2 _19347_ (
    .A(_8242_),
    .B(_8241_),
    .Y(_8243_)
);

FILL FILL_0__14197_ (
);

DFFSR _14482_ (
    .CLK(clk_bF$buf2),
    .D(_3672_[17]),
    .Q(\datapath_1.Data [17]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _14062_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3473_)
);

FILL FILL478040x182780 (
);

FILL FILL51680x266760 (
);

FILL FILL91200x375440 (
);

OR2X2 _15687_ (
    .A(_4637_),
    .B(_4636_),
    .Y(_4638_)
);

AND2X2 _15267_ (
    .A(_4202_),
    .B(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_4225_)
);

FILL FILL_1__17770_ (
);

FILL FILL_0__16763_ (
);

FILL FILL_0__16343_ (
);

FILL FILL74480x350740 (
);

FILL FILL492480x237120 (
);

DFFSR _8970_ (
    .CLK(clk_bF$buf32),
    .D(_201_[30]),
    .Q(\datapath_1.regfile_1.regOut[4] [30]),
    .R(rst_bF$buf93),
    .S(vdd)
);

OR2X2 _8550_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_65_)
);

OR2X2 _11187_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_1403_)
);

FILL FILL49400x143260 (
);

FILL FILL_1__13270_ (
);

FILL FILL_0__17968_ (
);

AND2X2 _17833_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_6752_)
);

OR2X2 _17413_ (
    .A(_6336_),
    .B(_6337_),
    .Y(_6338_)
);

FILL FILL_0__17128_ (
);

FILL FILL_0__12263_ (
);

AND2X2 _9755_ (
    .A(_668_),
    .B(_667_),
    .Y(_663_[2])
);

DFFSR _9335_ (
    .CLK(clk_bF$buf52),
    .D(_399_[8]),
    .Q(\datapath_1.regfile_1.regOut[7] [8]),
    .R(rst_bF$buf32),
    .S(vdd)
);

FILL FILL427120x340860 (
);

FILL FILL376960x59280 (
);

OR2X2 _18618_ (
    .A(_7524_),
    .B(_7521_),
    .Y(_7525_)
);

FILL FILL239400x172900 (
);

FILL FILL_0__13888_ (
);

FILL FILL_0__13468_ (
);

AND2X2 _13753_ (
    .A(_3084__bF$buf2),
    .B(\datapath_1.PCJump [23]),
    .Y(_3225_)
);

FILL FILL_0__13048_ (
);

OR2X2 _13333_ (
    .A(_2187_),
    .B(_2873_),
    .Y(_2874_)
);

FILL FILL_1__9497_ (
);

FILL FILL105640x79040 (
);

FILL FILL122360x29640 (
);

FILL FILL180880x113620 (
);

FILL FILL275120x251940 (
);

FILL FILL123120x158080 (
);

OR2X2 _14958_ (
    .A(\datapath_1.mux_pcsrc.dout [24]),
    .B(_4001__bF$buf3),
    .Y(_3985_)
);

OR2X2 _14538_ (
    .A(memoryOutData[13]),
    .B(_3803__bF$buf3),
    .Y(_3765_)
);

AND2X2 _14118_ (
    .A(_3352__bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3521_)
);

FILL FILL_1__16621_ (
);

FILL FILL503880x296400 (
);

FILL FILL_0__15614_ (
);

FILL FILL_1__19093_ (
);

AND2X2 _18791_ (
    .A(_6216__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_7695_)
);

FILL FILL_0__18086_ (
);

AND2X2 _18371_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_7282_)
);

FILL FILL283480x365560 (
);

DFFSR _10878_ (
    .CLK(clk_bF$buf71),
    .D(_1191_[3]),
    .Q(\datapath_1.regfile_1.regOut[19] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

OR2X2 _10458_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_1037_)
);

FILL FILL_1__17406_ (
);

OR2X2 _10038_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_817_)
);

FILL FILL_0__11954_ (
);

FILL FILL_0__11114_ (
);

FILL FILL15200x217360 (
);

OR2X2 _19156_ (
    .A(_8053_),
    .B(_8054_),
    .Y(_8055_)
);

FILL FILL126160x29640 (
);

OR2X2 _14291_ (
    .A(vdd),
    .B(ALUOut[17]),
    .Y(_3640_)
);

AND2X2 _8606_ (
    .A(_82_),
    .B(_81_),
    .Y(_69_[6])
);

FILL FILL41040x158080 (
);

FILL FILL253840x44460 (
);

FILL FILL_1__13746_ (
);

OR2X2 _12604_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2168_),
    .Y(_2169_)
);

FILL FILL381520x242060 (
);

FILL FILL230280x44460 (
);

FILL FILL428640x54340 (
);

OR2X2 _15496_ (
    .A(_4449_),
    .B(_4446_),
    .Y(_4450_)
);

AND2X2 _15076_ (
    .A(_4056_),
    .B(_4062_),
    .Y(_4063_)
);

FILL FILL_1__8768_ (
);

FILL FILL_0__16992_ (
);

FILL FILL_0__16572_ (
);

AND2X2 _13809_ (
    .A(_3084__bF$buf1),
    .B(\datapath_1.PCJump [31]),
    .Y(_3273_)
);

FILL FILL313880x266760 (
);

FILL FILL148200x197600 (
);

FILL FILL113240x83980 (
);

FILL FILL381520x108680 (
);

FILL FILL_0__17777_ (
);

FILL FILL194560x316160 (
);

OR2X2 _17642_ (
    .A(_6563_),
    .B(_6562_),
    .Y(_6564_)
);

FILL FILL_0__17357_ (
);

AND2X2 _17222_ (
    .A(_4208__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_6149_)
);

FILL FILL281960x321100 (
);

FILL FILL_0__12072_ (
);

DFFSR _9984_ (
    .CLK(clk_bF$buf28),
    .D(_729_[12]),
    .Q(\datapath_1.regfile_1.regOut[12] [12]),
    .R(rst_bF$buf96),
    .S(vdd)
);

OR2X2 _9564_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_581_)
);

OR2X2 _9144_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_361_)
);

FILL FILL277400x59280 (
);

FILL FILL_0__10805_ (
);

OR2X2 _18847_ (
    .A(_7746_),
    .B(_7749_),
    .Y(_7750_)
);

FILL FILL_0_BUFX2_insert641 (
);

INVX1 _18427_ (
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_7337_)
);

AND2X2 _18007_ (
    .A(_6232__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_6923_)
);

FILL FILL_0_BUFX2_insert643 (
);

AND2X2 _13982_ (
    .A(_3347__bF$buf0),
    .B(\datapath_1.PCJump [11]),
    .Y(_3404_)
);

FILL FILL_0__13697_ (
);

FILL FILL_0_BUFX2_insert645 (
);

FILL FILL_0__13277_ (
);

OR2X2 _13562_ (
    .A(ALUOut[24]),
    .B(_3079__bF$buf1),
    .Y(_3063_)
);

FILL FILL85120x360620 (
);

AOI21X1 _13142_ (
    .A(_2547_),
    .B(_2693_),
    .C(_2692_),
    .Y(_2694_)
);

FILL FILL_0_BUFX2_insert646 (
);

FILL FILL_0_BUFX2_insert647 (
);

FILL FILL120840x49400 (
);

FILL FILL_0_BUFX2_insert648 (
);

FILL FILL_0_BUFX2_insert649 (
);

FILL FILL399760x311220 (
);

FILL FILL_0__19503_ (
);

FILL FILL383800x197600 (
);

FILL FILL66120x197600 (
);

FILL FILL28120x79040 (
);

FILL FILL210520x256880 (
);

FILL FILL161120x301340 (
);

FILL FILL207480x207480 (
);

FILL FILL11400x247000 (
);

AND2X2 _14767_ (
    .A(_3877_),
    .B(_3876_),
    .Y(_3870_[3])
);

DFFSR _14347_ (
    .CLK(clk_bF$buf92),
    .D(_3606_[11]),
    .Q(ALUOut[11]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL_1__16010_ (
);

FILL FILL_0__15843_ (
);

AND2X2 _18180_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_7094_)
);

FILL FILL_1__17635_ (
);

OR2X2 _10687_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_1190__bF$buf0),
    .Y(_1150_)
);

OR2X2 _10267_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .B(_992__bF$buf2),
    .Y(_930_)
);

FILL FILL_0__16628_ (
);

AND2X2 _16913_ (
    .A(_4234__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_5845_)
);

FILL FILL_0__16208_ (
);

FILL FILL139080x93860 (
);

FILL FILL_0__11343_ (
);

AND2X2 _19385_ (
    .A(_6312__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_8280_)
);

FILL FILL209760x296400 (
);

DFFSR _8835_ (
    .CLK(clk_bF$buf97),
    .D(_135_[24]),
    .Q(\datapath_1.regfile_1.regOut[3] [24]),
    .R(rst_bF$buf77),
    .S(vdd)
);

BUFX2 _8415_ (
    .A(_1_[23]),
    .Y(memoryAddress[23])
);

FILL FILL329080x9880 (
);

FILL FILL_0__12968_ (
);

NAND3X1 _12833_ (
    .A(_2397_),
    .B(\datapath_1.alu_1.ALUInB [2]),
    .C(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2398_)
);

FILL FILL_0__12548_ (
);

AND2X2 _12413_ (
    .A(_2040_),
    .B(_2039_),
    .Y(_1983_[28])
);

FILL FILL455240x251940 (
);

FILL FILL420280x24700 (
);

FILL FILL_0__16381_ (
);

OR2X2 _13618_ (
    .A(_3109_),
    .B(_3106_),
    .Y(\datapath_1.mux_pcsrc.dout [3])
);

FILL FILL_1__18593_ (
);

OR2X2 _17871_ (
    .A(_6787_),
    .B(_6788_),
    .Y(_6789_)
);

FILL FILL_0__17586_ (
);

OR2X2 _17451_ (
    .A(_6374_),
    .B(_6375_),
    .Y(_6376_)
);

FILL FILL_0__17166_ (
);

OR2X2 _17031_ (
    .A(_5959_),
    .B(_5960_),
    .Y(_5961_)
);

FILL FILL367080x9880 (
);

FILL FILL275880x197600 (
);

OR2X2 _9793_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .B(_728__bF$buf1),
    .Y(_694_)
);

FILL FILL413440x113620 (
);

OR2X2 _9373_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .B(_530__bF$buf3),
    .Y(_474_)
);

FILL FILL_1__19378_ (
);

FILL FILL_0__10614_ (
);

FILL FILL424840x182780 (
);

AND2X2 _18656_ (
    .A(_6321__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_7562_)
);

AND2X2 _18236_ (
    .A(_6287__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_7149_)
);

AND2X2 _13791_ (
    .A(_3089__bF$buf1),
    .B(gnd),
    .Y(_3258_)
);

OR2X2 _13371_ (
    .A(_2908_),
    .B(_2376__bF$buf3),
    .Y(_2909_)
);

FILL FILL_0__9413_ (
);

FILL FILL_1__15298_ (
);

FILL FILL411160x187720 (
);

FILL FILL347320x360620 (
);

DFFSR _14996_ (
    .CLK(clk_bF$buf92),
    .D(_3936_[15]),
    .Q(\datapath_1.mux_iord.din0 [15]),
    .R(rst_bF$buf29),
    .S(vdd)
);

OR2X2 _14576_ (
    .A(IRWrite_bF$buf2),
    .B(\control_1.op [0]),
    .Y(_3790_)
);

OR2X2 _14156_ (
    .A(\datapath_1.Data [4]),
    .B(_3605__bF$buf1),
    .Y(_3549_)
);

FILL FILL_0__15232_ (
);

FILL FILL41800x296400 (
);

FILL FILL459800x276640 (
);

DFFSR _10496_ (
    .CLK(clk_bF$buf47),
    .D(_993_[8]),
    .Q(\datapath_1.regfile_1.regOut[16] [8]),
    .R(rst_bF$buf51),
    .S(vdd)
);

FILL FILL195320x271700 (
);

AND2X2 _10076_ (
    .A(_842_),
    .B(_841_),
    .Y(_795_[23])
);

FILL FILL_0__16857_ (
);

FILL FILL_0__16437_ (
);

AND2X2 _16722_ (
    .A(_4183__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_5657_)
);

OR2X2 _16302_ (
    .A(_5242_),
    .B(_5243_),
    .Y(_5244_)
);

FILL FILL_0__11992_ (
);

OR2X2 _19194_ (
    .A(_8091_),
    .B(_8078_),
    .Y(_8092_)
);

OR2X2 _8644_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .B(_134__bF$buf0),
    .Y(_108_)
);

FILL FILL_1__13364_ (
);

OR2X2 _17927_ (
    .A(_6844_),
    .B(_6829_),
    .Y(_6845_)
);

AND2X2 _17507_ (
    .A(_6259__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_6431_)
);

OR2X2 _12642_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2206_),
    .Y(_2207_)
);

FILL FILL_0__12357_ (
);

OR2X2 _12222_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_1933_)
);

FILL FILL230280x182780 (
);

DFFSR _9849_ (
    .CLK(clk_bF$buf36),
    .D(_663_[6]),
    .Q(\datapath_1.regfile_1.regOut[11] [6]),
    .R(rst_bF$buf25),
    .S(vdd)
);

OR2X2 _9429_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_511_)
);

OR2X2 _9009_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_291_)
);

FILL FILL_0__16190_ (
);

FILL FILL_1__14569_ (
);

FILL FILL303240x296400 (
);

OR2X2 _13847_ (
    .A(\datapath_1.a [10]),
    .B(_3342__bF$buf2),
    .Y(_3298_)
);

AND2X2 _13427_ (
    .A(_2961_),
    .B(_2958_),
    .Y(_2962_)
);

NOR2X1 _13007_ (
    .A(_2566_),
    .B(_2564_),
    .Y(_2567_)
);

FILL FILL_0__14923_ (
);

FILL FILL_0__14503_ (
);

FILL FILL114000x98800 (
);

OR2X2 _17680_ (
    .A(_6599_),
    .B(_6600_),
    .Y(_6601_)
);

AND2X2 _17260_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_6187_)
);

FILL FILL284240x118560 (
);

FILL FILL371640x123500 (
);

AND2X2 _9182_ (
    .A(_386_),
    .B(_385_),
    .Y(_333_[26])
);

FILL FILL_1__11430_ (
);

FILL FILL_0__15708_ (
);

FILL FILL_0__10423_ (
);

OR2X2 _18885_ (
    .A(_7780_),
    .B(_7787_),
    .Y(_7788_)
);

OR2X2 _18465_ (
    .A(_7373_),
    .B(_7366_),
    .Y(_7374_)
);

AND2X2 _18045_ (
    .A(_6229__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_6961_)
);

FILL FILL438520x296400 (
);

OR2X2 _13180_ (
    .A(_2224_),
    .B(_2210_),
    .Y(_2729_)
);

FILL FILL_0__19121_ (
);

FILL FILL47880x365560 (
);

FILL FILL_0__11628_ (
);

DFFSR _11913_ (
    .CLK(clk_bF$buf49),
    .D(_1719_[6]),
    .Q(\datapath_1.regfile_1.regOut[27] [6]),
    .R(rst_bF$buf106),
    .S(vdd)
);

OR2X2 _14385_ (
    .A(memoryOutData[5]),
    .B(_3737__bF$buf1),
    .Y(_3683_)
);

FILL FILL_0__15881_ (
);

FILL FILL_0__15461_ (
);

FILL FILL10640x108680 (
);

FILL FILL200640x271700 (
);

FILL FILL276640x133380 (
);

FILL FILL_0__16666_ (
);

OR2X2 _16951_ (
    .A(_5875_),
    .B(_5882_),
    .Y(_5883_)
);

OR2X2 _16531_ (
    .A(_5468_),
    .B(_5467_),
    .Y(_5469_)
);

FILL FILL_0__16246_ (
);

OR2X2 _16111_ (
    .A(_5055_),
    .B(_5052_),
    .Y(_5056_)
);

FILL FILL449920x153140 (
);

AND2X2 _8873_ (
    .A(_220_),
    .B(_219_),
    .Y(_201_[9])
);

BUFX2 _8453_ (
    .A(_2_[29]),
    .Y(memoryWriteData[29])
);

FILL FILL349600x247000 (
);

FILL FILL_1__18458_ (
);

FILL FILL306280x79040 (
);

AND2X2 _17736_ (
    .A(_6211__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_6656_)
);

OR2X2 _17316_ (
    .A(_6241_),
    .B(_6224_),
    .Y(_6242_)
);

FILL FILL18240x271700 (
);

FILL FILL31920x44460 (
);

OR2X2 _12871_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2436_)
);

DFFSR _12451_ (
    .CLK(clk_bF$buf72),
    .D(_1983_[28]),
    .Q(\datapath_1.regfile_1.regOut[31] [28]),
    .R(rst_bF$buf32),
    .S(vdd)
);

OR2X2 _12031_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .B(_1850__bF$buf2),
    .Y(_1846_)
);

FILL FILL383800x98800 (
);

OR2X2 _9658_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .B(_662__bF$buf3),
    .Y(_624_)
);

OR2X2 _9238_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .B(_464__bF$buf3),
    .Y(_404_)
);

FILL FILL_1__11906_ (
);

FILL FILL_1__14378_ (
);

OR2X2 _13656_ (
    .A(_3140_),
    .B(_3141_),
    .Y(_3142_)
);

MUX2X1 _13236_ (
    .A(_2501_),
    .B(_2376__bF$buf0),
    .S(_2781_),
    .Y(_2782_)
);

FILL FILL_0__14312_ (
);

FILL FILL19000x69160 (
);

FILL FILL380760x0 (
);

FILL FILL_1__16104_ (
);

FILL FILL98040x148200 (
);

FILL FILL_0__15937_ (
);

AND2X2 _15802_ (
    .A(_4751_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [8])
);

FILL FILL_0__10652_ (
);

FILL FILL242440x207480 (
);

OR2X2 _18694_ (
    .A(_7599_),
    .B(_7598_),
    .Y(_7600_)
);

OR2X2 _18274_ (
    .A(_7184_),
    .B(_7185_),
    .Y(_7186_)
);

FILL FILL_0__19350_ (
);

FILL FILL_1__12864_ (
);

FILL FILL_1__12024_ (
);

FILL FILL185440x158080 (
);

FILL FILL_0__11857_ (
);

FILL FILL_0__9451_ (
);

OR2X2 _11722_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .B(_1718__bF$buf2),
    .Y(_1680_)
);

FILL FILL_0__11437_ (
);

OR2X2 _11302_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .B(_1520__bF$buf2),
    .Y(_1460_)
);

FILL FILL310080x276640 (
);

OR2X2 _19479_ (
    .A(gnd),
    .B(_8385__bF$buf0),
    .Y(_8355_)
);

OR2X2 _19059_ (
    .A(_7957_),
    .B(_7958_),
    .Y(_7959_)
);

OR2X2 _14194_ (
    .A(MemToReg_bF$buf3),
    .B(ALUOut[17]),
    .Y(_3574_)
);

OR2X2 _8929_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_266__bF$buf4),
    .Y(_258_)
);

OR2X2 _8509_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .B(_68__bF$buf4),
    .Y(_38_)
);

FILL FILL227240x286520 (
);

FILL FILL_0__15690_ (
);

FILL FILL_1_BUFX2_insert570 (
);

XNOR2X1 _12927_ (
    .A(_2160_),
    .B(_2491_),
    .Y(_2492_)
);

FILL FILL244720x296400 (
);

NOR2X1 _12507_ (
    .A(\control_1.reg_state.dout [1]),
    .B(\control_1.reg_state.dout [0]),
    .Y(_2103_)
);

FILL FILL10640x24700 (
);

FILL FILL_1_BUFX2_insert578 (
);

OR2X2 _15399_ (
    .A(_4354_),
    .B(_4351_),
    .Y(_4355_)
);

FILL FILL490960x153140 (
);

FILL FILL_0__16895_ (
);

OR2X2 _16760_ (
    .A(_5694_),
    .B(_5679_),
    .Y(_5695_)
);

FILL FILL_0__16055_ (
);

AND2X2 _16340_ (
    .A(_4175__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_5281_)
);

DFFSR _8682_ (
    .CLK(clk_bF$buf19),
    .D(_69_[0]),
    .Q(\datapath_1.regfile_1.regOut[2] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

BUFX2 BUFX2_insert240 (
    .A(_6236_),
    .Y(_6236__bF$buf3)
);

BUFX2 BUFX2_insert241 (
    .A(_6236_),
    .Y(_6236__bF$buf2)
);

BUFX2 BUFX2_insert242 (
    .A(_6236_),
    .Y(_6236__bF$buf1)
);

BUFX2 BUFX2_insert243 (
    .A(_6236_),
    .Y(_6236__bF$buf0)
);

BUFX2 BUFX2_insert244 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf4 )
);

AND2X2 _17965_ (
    .A(_6289__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_6882_)
);

FILL FILL134520x316160 (
);

AND2X2 _17545_ (
    .A(_6211__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_6468_)
);

BUFX2 BUFX2_insert245 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf3 )
);

BUFX2 BUFX2_insert246 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf2 )
);

AND2X2 _17125_ (
    .A(_4135__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_6054_)
);

FILL FILL221920x321100 (
);

BUFX2 BUFX2_insert247 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf1 )
);

BUFX2 BUFX2_insert248 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf0 )
);

FILL FILL_0__12395_ (
);

OR2X2 _12680_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(_2244_),
    .Y(_2245_)
);

BUFX2 BUFX2_insert249 (
    .A(_4146_),
    .Y(_4146__bF$buf4)
);

AND2X2 _12260_ (
    .A(_1958_),
    .B(_1957_),
    .Y(_1917_[20])
);

FILL FILL_0__18621_ (
);

FILL FILL438520x14820 (
);

FILL FILL_0__18201_ (
);

AND2X2 _9887_ (
    .A(_736_),
    .B(_735_),
    .Y(_729_[3])
);

DFFSR _9467_ (
    .CLK(clk_bF$buf57),
    .D(_465_[11]),
    .Q(\datapath_1.regfile_1.regOut[8] [11]),
    .R(rst_bF$buf81),
    .S(vdd)
);

AND2X2 _9047_ (
    .A(_316_),
    .B(_315_),
    .Y(_267_[24])
);

FILL FILL_1__11715_ (
);

FILL FILL_0__10708_ (
);

FILL FILL_1__14187_ (
);

OR2X2 _13885_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [23]),
    .Y(_3323_)
);

AND2X2 _13465_ (
    .A(_2997_),
    .B(_2994_),
    .Y(_2998_)
);

OR2X2 _13045_ (
    .A(_2275_),
    .B(_2601_),
    .Y(_2602_)
);

FILL FILL_0__19406_ (
);

FILL FILL_0__14961_ (
);

FILL FILL_0__14541_ (
);

FILL FILL98800x335920 (
);

FILL FILL_0__14121_ (
);

FILL FILL238640x330980 (
);

FILL FILL_0__9507_ (
);

FILL FILL183160x207480 (
);

FILL FILL_1__16753_ (
);

FILL FILL208240x88920 (
);

FILL FILL356440x227240 (
);

FILL FILL_0__15746_ (
);

FILL FILL_0__15326_ (
);

AND2X2 _15611_ (
    .A(_4160__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_4563_)
);

FILL FILL_0__10041_ (
);

FILL FILL342760x251940 (
);

AND2X2 _18083_ (
    .A(_6297__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_6998_)
);

FILL FILL443080x138320 (
);

FILL FILL_1__17958_ (
);

AND2X2 _16816_ (
    .A(_4234__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_5750_)
);

FILL FILL73720x247000 (
);

FILL FILL396720x321100 (
);

FILL FILL_0__9680_ (
);

AND2X2 _11951_ (
    .A(_1792_),
    .B(_1791_),
    .Y(_1785_[3])
);

DFFSR _11531_ (
    .CLK(clk_bF$buf82),
    .D(_1521_[11]),
    .Q(\datapath_1.regfile_1.regOut[24] [11]),
    .R(rst_bF$buf39),
    .S(vdd)
);

FILL FILL_0__11246_ (
);

AND2X2 _11111_ (
    .A(_1372_),
    .B(_1371_),
    .Y(_1323_[24])
);

AND2X2 _19288_ (
    .A(_6238__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_8185_)
);

AND2X2 _8738_ (
    .A(_150_),
    .B(_149_),
    .Y(_135_[7])
);

FILL FILL323000x212420 (
);

FILL FILL_1__13038_ (
);

AND2X2 _12736_ (
    .A(_2298_),
    .B(_2300_),
    .Y(_2301_)
);

DFFSR _12316_ (
    .CLK(clk_bF$buf110),
    .D(_1917_[22]),
    .Q(\datapath_1.regfile_1.regOut[30] [22]),
    .R(rst_bF$buf50),
    .S(vdd)
);

FILL FILL300960x113620 (
);

FILL FILL141360x93860 (
);

FILL FILL_0__13812_ (
);

FILL FILL269040x79040 (
);

FILL FILL_0__16284_ (
);

FILL FILL348840x242060 (
);

FILL FILL242440x4940 (
);

FILL FILL_1__9001_ (
);

FILL FILL285760x54340 (
);

OR2X2 _8491_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .B(_68__bF$buf0),
    .Y(_26_)
);

FILL FILL_1__15604_ (
);

FILL FILL_1__18076_ (
);

FILL FILL179360x143260 (
);

FILL FILL147440x355680 (
);

AND2X2 _17774_ (
    .A(_6302__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_6694_)
);

FILL FILL_0__17069_ (
);

AND2X2 _17354_ (
    .A(_6279_),
    .B(_6278_),
    .Y(_6280_)
);

FILL FILL_0__18850_ (
);

FILL FILL_0__18010_ (
);

OR2X2 _9696_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_649_)
);

OR2X2 _9276_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_429_)
);

FILL FILL_0__10937_ (
);

AND2X2 _10802_ (
    .A(_1206_),
    .B(_1205_),
    .Y(_1191_[7])
);

AND2X2 _18979_ (
    .A(_6232__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [25]),
    .Y(_7880_)
);

OR2X2 _18559_ (
    .A(_7466_),
    .B(_7465_),
    .Y(_7467_)
);

OR2X2 _18139_ (
    .A(_7049_),
    .B(_7052_),
    .Y(_7053_)
);

OR2X2 _13694_ (
    .A(_3174_),
    .B(_3173_),
    .Y(_3175_)
);

AND2X2 _13274_ (
    .A(_2817_),
    .B(_2815_),
    .Y(_2818_)
);

FILL FILL_0__19215_ (
);

OR2X2 _19500_ (
    .A(gnd),
    .B(_8385__bF$buf0),
    .Y(_8369_)
);

FILL FILL_0__14770_ (
);

FILL FILL_1__12729_ (
);

FILL FILL353400x64220 (
);

FILL FILL_0__9316_ (
);

FILL FILL332120x143260 (
);

AND2X2 _14899_ (
    .A(_3945_),
    .B(_3944_),
    .Y(_3936_[4])
);

DFFSR _14479_ (
    .CLK(clk_bF$buf65),
    .D(_3672_[14]),
    .Q(\datapath_1.Data [14]),
    .R(rst_bF$buf36),
    .S(vdd)
);

AND2X2 _14059_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3470_)
);

FILL FILL69920x370500 (
);

FILL FILL_0__15975_ (
);

FILL FILL501600x108680 (
);

OR2X2 _15840_ (
    .A(_4785_),
    .B(_4788_),
    .Y(_4789_)
);

FILL FILL_0__15555_ (
);

AND2X2 _15420_ (
    .A(_4158__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_4375_)
);

FILL FILL82840x365560 (
);

DFFSR _15000_ (
    .CLK(clk_bF$buf77),
    .D(_3936_[19]),
    .Q(\datapath_1.mux_iord.din0 [19]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL_0__10690_ (
);

FILL FILL314640x316160 (
);

FILL FILL304000x276640 (
);

FILL FILL456000x0 (
);

OR2X2 _10399_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .B(_1058__bF$buf0),
    .Y(_998_)
);

FILL FILL_1__12482_ (
);

AND2X2 _16625_ (
    .A(_4210__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_5562_)
);

AND2X2 _16205_ (
    .A(_4160__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_5148_)
);

FILL FILL145160x217360 (
);

OR2X2 _11760_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_1705_)
);

FILL FILL_0__11475_ (
);

OR2X2 _11340_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_1485_)
);

FILL FILL_0__11055_ (
);

OR2X2 _19097_ (
    .A(_7981_),
    .B(_7996_),
    .Y(_7997_)
);

FILL FILL23560x217360 (
);

DFFSR _8967_ (
    .CLK(clk_bF$buf49),
    .D(_201_[27]),
    .Q(\datapath_1.regfile_1.regOut[4] [27]),
    .R(rst_bF$buf106),
    .S(vdd)
);

OR2X2 _8547_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_63_)
);

FILL FILL87400x93860 (
);

FILL FILL327560x128440 (
);

FILL FILL_1__13687_ (
);

FILL FILL418760x330980 (
);

FILL FILL_1_BUFX2_insert950 (
);

AND2X2 _12965_ (
    .A(_2527_),
    .B(_2515_),
    .Y(_2528_)
);

NOR3X1 _12545_ (
    .A(_2113_),
    .B(_2133_),
    .C(_2132_),
    .Y(_2134_)
);

AND2X2 _12125_ (
    .A(_1888_),
    .B(_1887_),
    .Y(_1851_[18])
);

FILL FILL_1_BUFX2_insert958 (
);

FILL FILL_0__18906_ (
);

FILL FILL_0__13201_ (
);

FILL FILL490200x321100 (
);

FILL FILL380760x217360 (
);

BUFX2 BUFX2_insert620 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf19)
);

BUFX2 BUFX2_insert621 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf18)
);

BUFX2 BUFX2_insert622 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf17)
);

BUFX2 BUFX2_insert623 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf16)
);

BUFX2 BUFX2_insert624 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf15)
);

AND2X2 _17583_ (
    .A(_6264__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_6506_)
);

BUFX2 BUFX2_insert625 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf14)
);

FILL FILL_0__17298_ (
);

BUFX2 BUFX2_insert626 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf13)
);

AND2X2 _17163_ (
    .A(_4223__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_6091_)
);

BUFX2 BUFX2_insert627 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf12)
);

BUFX2 BUFX2_insert628 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf11)
);

BUFX2 BUFX2_insert629 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf10)
);

FILL FILL348080x286520 (
);

FILL FILL110200x370500 (
);

FILL FILL101840x247000 (
);

FILL FILL142880x34580 (
);

FILL FILL192280x276640 (
);

FILL FILL120080x316160 (
);

DFFSR _9085_ (
    .CLK(clk_bF$buf5),
    .D(_267_[16]),
    .Q(\datapath_1.regfile_1.regOut[5] [16]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL_1__11333_ (
);

FILL FILL365560x296400 (
);

FILL FILL15960x232180 (
);

FILL FILL_0__8760_ (
);

FILL FILL_0__10326_ (
);

OR2X2 _10611_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_1119_)
);

FILL FILL503120x212420 (
);

OR2X2 _18788_ (
    .A(_7691_),
    .B(_7690_),
    .Y(_7692_)
);

AND2X2 _18368_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_7279_)
);

FILL FILL247000x202540 (
);

XOR2X1 _13083_ (
    .A(_2269_),
    .B(_2637_),
    .Y(_2638_)
);

FILL FILL_0__19444_ (
);

FILL FILL224960x103740 (
);

FILL FILL414200x375440 (
);

AND2X2 _11816_ (
    .A(_1722_),
    .B(_1721_),
    .Y(_1719_[1])
);

FILL FILL_0__9125_ (
);

OR2X2 _14288_ (
    .A(vdd),
    .B(ALUOut[16]),
    .Y(_3638_)
);

FILL FILL_0__15784_ (
);

FILL FILL_0__15364_ (
);

FILL FILL272840x326040 (
);

FILL FILL_1__17576_ (
);

OR2X2 _16854_ (
    .A(_5785_),
    .B(_5786_),
    .Y(_5787_)
);

OR2X2 _16434_ (
    .A(_5372_),
    .B(_5373_),
    .Y(_5374_)
);

FILL FILL_0__16149_ (
);

AND2X2 _16014_ (
    .A(_4135__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_4960_)
);

FILL FILL_0__17510_ (
);

FILL FILL36480x256880 (
);

OR2X2 _8776_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .B(_200__bF$buf2),
    .Y(_176_)
);

FILL FILL382280x321100 (
);

FILL FILL_1__10604_ (
);

FILL FILL427880x172900 (
);

OR2X2 _17639_ (
    .A(_6559_),
    .B(_6560_),
    .Y(_6561_)
);

AND2X2 _17219_ (
    .A(_4197__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_6146_)
);

NAND3X1 _12774_ (
    .A(_2330_),
    .B(\datapath_1.alu_1.ALUInA [24]),
    .C(_2333_),
    .Y(_2339_)
);

FILL FILL_0__12489_ (
);

OR2X2 _12354_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_2001_)
);

FILL FILL477280x227240 (
);

FILL FILL357960x177840 (
);

FILL FILL_0__18715_ (
);

FILL FILL_0__13850_ (
);

FILL FILL_0__13430_ (
);

FILL FILL76760x350740 (
);

FILL FILL503880x24700 (
);

FILL FILL308560x301340 (
);

OR2X2 _13979_ (
    .A(_3401_),
    .B(_3400_),
    .Y(_3402_)
);

OR2X2 _13559_ (
    .A(ALUOut[23]),
    .B(_3079__bF$buf4),
    .Y(_3061_)
);

AOI22X1 _13139_ (
    .A(_2690_),
    .B(_2379__bF$buf0),
    .C(_2593_),
    .D(_2687_),
    .Y(_2691_)
);

FILL FILL_1__15222_ (
);

AND2X2 _14920_ (
    .A(_3959_),
    .B(_3958_),
    .Y(_3936_[11])
);

AND2X2 _14500_ (
    .A(_3739_),
    .B(_3802_),
    .Y(_3738_[0])
);

FILL FILL250800x34580 (
);

AND2X2 _17392_ (
    .A(_6317__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_6318_)
);

FILL FILL503880x207480 (
);

FILL FILL429400x340860 (
);

FILL FILL_1__16427_ (
);

FILL FILL273600x330980 (
);

OR2X2 _15705_ (
    .A(_4640_),
    .B(_4655_),
    .Y(_4656_)
);

FILL FILL_0__10975_ (
);

OR2X2 _10840_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .B(_1256__bF$buf3),
    .Y(_1232_)
);

FILL FILL_0__10555_ (
);

FILL FILL137560x370500 (
);

OR2X2 _10420_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .B(_1058__bF$buf0),
    .Y(_1012_)
);

FILL FILL_0__10135_ (
);

FILL FILL254600x167960 (
);

DFFSR _10000_ (
    .CLK(clk_bF$buf72),
    .D(_729_[28]),
    .Q(\datapath_1.regfile_1.regOut[12] [28]),
    .R(rst_bF$buf32),
    .S(vdd)
);

INVX1 _18597_ (
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_7504_)
);

FILL FILL24320x172900 (
);

OR2X2 _18177_ (
    .A(_7087_),
    .B(_7090_),
    .Y(_7091_)
);

FILL FILL351880x118560 (
);

OR2X2 _11625_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_1635_)
);

OR2X2 _11205_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_1415_)
);

FILL FILL111720x182780 (
);

AND2X2 _14097_ (
    .A(_3352__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3503_)
);

FILL FILL_0__12701_ (
);

FILL FILL_1__16180_ (
);

FILL FILL32680x286520 (
);

FILL FILL_0__15173_ (
);

FILL FILL285760x365560 (
);

FILL FILL180880x187720 (
);

FILL FILL424080x54340 (
);

FILL FILL_0__16798_ (
);

OR2X2 _16663_ (
    .A(_5595_),
    .B(_5598_),
    .Y(_5599_)
);

FILL FILL_0__16378_ (
);

AND2X2 _16243_ (
    .A(_4223__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_5186_)
);

FILL FILL131480x311220 (
);

FILL FILL_0__11093_ (
);

OR2X2 _8585_ (
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .Y(_133_)
);

FILL FILL_1__10413_ (
);

FILL FILL383800x242060 (
);

OR2X2 _17868_ (
    .A(_6784_),
    .B(_6785_),
    .Y(_6786_)
);

FILL FILL253080x44460 (
);

OR2X2 _17448_ (
    .A(_6369_),
    .B(_6372_),
    .Y(_6373_)
);

OR2X2 _17028_ (
    .A(_5956_),
    .B(_5957_),
    .Y(_5958_)
);

AND2X2 _12583_ (
    .A(_2152_),
    .B(_2151_),
    .Y(_2143_[3])
);

OR2X2 _12163_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .B(_1916__bF$buf0),
    .Y(_1914_)
);

FILL FILL_0__18944_ (
);

FILL FILL44080x14820 (
);

FILL FILL_0__18524_ (
);

FILL FILL343520x83980 (
);

FILL FILL_1__11618_ (
);

FILL FILL383800x108680 (
);

FILL FILL250800x197600 (
);

AND2X2 _13788_ (
    .A(_3084__bF$buf1),
    .B(\datapath_1.PCJump [28]),
    .Y(_3255_)
);

FILL FILL256120x271700 (
);

XOR2X1 _13368_ (
    .A(_2402_),
    .B(_2185_),
    .Y(_2906_)
);

FILL FILL_1__15871_ (
);

FILL FILL_0__19309_ (
);

FILL FILL196840x316160 (
);

FILL FILL_0__14444_ (
);

FILL FILL_0__14024_ (
);

FILL FILL440800x14820 (
);

CLKBUF1 CLKBUF1_insert160 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf63)
);

CLKBUF1 CLKBUF1_insert161 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf62)
);

CLKBUF1 CLKBUF1_insert162 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf61)
);

CLKBUF1 CLKBUF1_insert163 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf60)
);

FILL FILL21280x88920 (
);

CLKBUF1 CLKBUF1_insert164 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf59)
);

CLKBUF1 CLKBUF1_insert165 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf58)
);

CLKBUF1 CLKBUF1_insert166 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert167 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert168 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf55)
);

FILL FILL283480x227240 (
);

CLKBUF1 CLKBUF1_insert169 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf54)
);

FILL FILL493240x103740 (
);

AND2X2 _15934_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_4881_)
);

FILL FILL_0__15649_ (
);

FILL FILL347320x83980 (
);

AND2X2 _15514_ (
    .A(_4200__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_4468_)
);

FILL FILL_0__15229_ (
);

FILL FILL87400x360620 (
);

FILL FILL_0__10784_ (
);

FILL FILL68400x197600 (
);

FILL FILL_0__19482_ (
);

FILL FILL_0__19062_ (
);

FILL FILL505400x326040 (
);

FILL FILL_1__12576_ (
);

OR2X2 _16719_ (
    .A(_5652_),
    .B(_5653_),
    .Y(_5654_)
);

FILL FILL_0__9583_ (
);

FILL FILL_0__11989_ (
);

OR2X2 _11854_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .B(_1784__bF$buf3),
    .Y(_1748_)
);

FILL FILL_0__9163_ (
);

FILL FILL_0__11569_ (
);

OR2X2 _11434_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .B(_1586__bF$buf2),
    .Y(_1528_)
);

DFFSR _11014_ (
    .CLK(clk_bF$buf107),
    .D(_1257_[10]),
    .Q(\datapath_1.regfile_1.regOut[20] [10]),
    .R(rst_bF$buf37),
    .S(vdd)
);

FILL FILL_0__12930_ (
);

FILL FILL_0__12510_ (
);

FILL FILL127680x113620 (
);

FILL FILL82080x79040 (
);

FILL FILL108680x271700 (
);

OR2X2 _12639_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(_2203_),
    .Y(_2204_)
);

FILL FILL178600x291460 (
);

OR2X2 _12219_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_1931_)
);

FILL FILL_1__14722_ (
);

FILL FILL467400x306280 (
);

FILL FILL_0__13715_ (
);

FILL FILL_1__17194_ (
);

FILL FILL302480x9880 (
);

AND2X2 _16892_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_5824_)
);

OR2X2 _16472_ (
    .A(_5403_),
    .B(_5410_),
    .Y(_5411_)
);

FILL FILL_0__16187_ (
);

AND2X2 _16052_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_4998_)
);

FILL FILL62320x138320 (
);

FILL FILL361000x44460 (
);

BUFX2 _8394_ (
    .A(_1_[2]),
    .Y(memoryAddress[2])
);

FILL FILL_1__18399_ (
);

FILL FILL79040x281580 (
);

FILL FILL142880x197600 (
);

OR2X2 _17677_ (
    .A(_6594_),
    .B(_6597_),
    .Y(_6598_)
);

AND2X2 _17257_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_6184_)
);

AND2X2 _12392_ (
    .A(_2026_),
    .B(_2025_),
    .Y(_1983_[21])
);

FILL FILL_1__19340_ (
);

FILL FILL62320x49400 (
);

FILL FILL_0__18333_ (
);

DFFSR _9599_ (
    .CLK(clk_bF$buf22),
    .D(_531_[14]),
    .Q(\datapath_1.regfile_1.regOut[9] [14]),
    .R(rst_bF$buf7),
    .S(vdd)
);

AND2X2 _9179_ (
    .A(_384_),
    .B(_383_),
    .Y(_333_[25])
);

FILL FILL_0__8854_ (
);

FILL FILL_0__8434_ (
);

OR2X2 _10705_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .B(_1190__bF$buf0),
    .Y(_1162_)
);

FILL FILL383040x286520 (
);

FILL FILL_0_BUFX2_insert990 (
);

FILL FILL_0_BUFX2_insert991 (
);

FILL FILL_0_BUFX2_insert992 (
);

FILL FILL_0_BUFX2_insert993 (
);

OR2X2 _13597_ (
    .A(_3091_),
    .B(_3086_),
    .Y(\datapath_1.mux_pcsrc.dout [0])
);

FILL FILL_0_BUFX2_insert995 (
);

AND2X2 _13177_ (
    .A(_2726_),
    .B(_2716_),
    .Y(_2727_)
);

FILL FILL_0_BUFX2_insert997 (
);

FILL FILL_0_BUFX2_insert999 (
);

AND2X2 _19403_ (
    .A(_6238__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_8298_)
);

FILL FILL_0__14673_ (
);

FILL FILL50920x232180 (
);

FILL FILL_0__14253_ (
);

FILL FILL_0__9639_ (
);

FILL FILL_1__16045_ (
);

FILL FILL309320x266760 (
);

FILL FILL_0__15878_ (
);

AND2X2 _15743_ (
    .A(_4197__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_4693_)
);

AND2X2 _15323_ (
    .A(_4175__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_4280_)
);

FILL FILL_0__15038_ (
);

FILL FILL_0__10173_ (
);

FILL FILL_0__19291_ (
);

FILL FILL176320x340860 (
);

FILL FILL_1__12385_ (
);

AND2X2 _16948_ (
    .A(_4130__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_5880_)
);

OR2X2 _16528_ (
    .A(_5462_),
    .B(_5465_),
    .Y(_5466_)
);

AND2X2 _16108_ (
    .A(_4187__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_5053_)
);

DFFSR _11663_ (
    .CLK(clk_bF$buf67),
    .D(_1587_[14]),
    .Q(\datapath_1.regfile_1.regOut[25] [14]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL_0__11378_ (
);

AND2X2 _11243_ (
    .A(_1440_),
    .B(_1439_),
    .Y(_1389_[25])
);

FILL FILL_0__17604_ (
);

FILL FILL193040x256880 (
);

OR2X2 _9811_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .B(_728__bF$buf3),
    .Y(_706_)
);

OR2X2 _12868_ (
    .A(_2431_),
    .B(_2432_),
    .Y(_2433_)
);

DFFSR _12448_ (
    .CLK(clk_bF$buf69),
    .D(_1983_[25]),
    .Q(\datapath_1.regfile_1.regOut[31] [25]),
    .R(rst_bF$buf79),
    .S(vdd)
);

OR2X2 _12028_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .B(_1850__bF$buf0),
    .Y(_1844_)
);

FILL FILL_1__14531_ (
);

FILL FILL_0__18809_ (
);

FILL FILL_0__13944_ (
);

FILL FILL_0__13524_ (
);

FILL FILL375440x167960 (
);

FILL FILL_0__13104_ (
);

OR2X2 _16281_ (
    .A(_5207_),
    .B(_5222_),
    .Y(_5223_)
);

FILL FILL_1__9133_ (
);

INVX1 _17486_ (
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_6410_)
);

FILL FILL106400x335920 (
);

AND2X2 _17066_ (
    .A(_4146__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_5996_)
);

FILL FILL_0__18982_ (
);

FILL FILL_0__18562_ (
);

AND2X2 _10934_ (
    .A(_1274_),
    .B(_1273_),
    .Y(_1257_[8])
);

DFFSR _10514_ (
    .CLK(clk_bF$buf109),
    .D(_993_[26]),
    .Q(\datapath_1.regfile_1.regOut[16] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL209000x34580 (
);

FILL FILL356440x113620 (
);

FILL FILL_0__19347_ (
);

INVX1 _19212_ (
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_8110_)
);

FILL FILL367840x182780 (
);

FILL FILL286520x118560 (
);

FILL FILL_0__9448_ (
);

FILL FILL_0__9028_ (
);

OR2X2 _11719_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .B(_1718__bF$buf3),
    .Y(_1678_)
);

FILL FILL373920x123500 (
);

FILL FILL24320x335920 (
);

FILL FILL_1__16694_ (
);

AND2X2 _15972_ (
    .A(_4154__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_4919_)
);

FILL FILL_0__15267_ (
);

OR2X2 _15552_ (
    .A(_4503_),
    .B(_4504_),
    .Y(_4505_)
);

NOR2X1 _15132_ (
    .A(_4033_),
    .B(_4065__bF$buf2),
    .Y(\datapath_1.regfile_1.regEn [16])
);

FILL FILL305520x9880 (
);

FILL FILL_1__17059_ (
);

OR2X2 _16757_ (
    .A(_5690_),
    .B(_5691_),
    .Y(_5692_)
);

AND2X2 _16337_ (
    .A(_4230__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_5278_)
);

OR2X2 _11892_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_1773_)
);

FILL FILL_0__11187_ (
);

OR2X2 _11472_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_1553_)
);

OR2X2 _11052_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_1333_)
);

FILL FILL_0__17833_ (
);

FILL FILL_0__17413_ (
);

OR2X2 _8679_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_131_)
);

FILL FILL322240x321100 (
);

AND2X2 _9620_ (
    .A(_598_),
    .B(_661_),
    .Y(_597_[0])
);

DFFSR _9200_ (
    .CLK(clk_bF$buf17),
    .D(_333_[2]),
    .Q(\datapath_1.regfile_1.regOut[6] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _12677_ (
    .A(_2234_),
    .B(_2241_),
    .Y(_2242_)
);

FILL FILL_1__19205_ (
);

AND2X2 _12257_ (
    .A(_1956_),
    .B(_1955_),
    .Y(_1917_[19])
);

OR2X2 _18903_ (
    .A(_7773_),
    .B(_7805_),
    .Y(_7806_)
);

FILL FILL_0__13753_ (
);

AND2X2 _16090_ (
    .A(_4158__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_5035_)
);

FILL FILL_0__8719_ (
);

FILL FILL478800x34580 (
);

FILL FILL_1__15545_ (
);

FILL FILL457520x321100 (
);

OR2X2 _14823_ (
    .A(\datapath_1.rd2 [22]),
    .B(_3935__bF$buf4),
    .Y(_3915_)
);

FILL FILL_0__14538_ (
);

FILL FILL_0__14118_ (
);

OR2X2 _14403_ (
    .A(memoryOutData[11]),
    .B(_3737__bF$buf0),
    .Y(_3695_)
);

AND2X2 _17295_ (
    .A(_6220_),
    .B(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_6221_)
);

FILL FILL282720x148200 (
);

FILL FILL288040x222300 (
);

FILL FILL383040x98800 (
);

FILL FILL_1__11465_ (
);

OR2X2 _15608_ (
    .A(_4545_),
    .B(_4560_),
    .Y(_4561_)
);

FILL FILL_0__8892_ (
);

FILL FILL_0__10458_ (
);

OR2X2 _10743_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_1187_)
);

OR2X2 _10323_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_967_)
);

FILL FILL468920x256880 (
);

AND2X2 _19441_ (
    .A(_8329_),
    .B(_8328_),
    .Y(_8320_[4])
);

FILL FILL_0__19156_ (
);

AND2X2 _19021_ (
    .A(_6317__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_7922_)
);

FILL FILL_0__14291_ (
);

FILL FILL_0__9257_ (
);

AND2X2 _11948_ (
    .A(_1790_),
    .B(_1789_),
    .Y(_1785_[2])
);

DFFSR _11528_ (
    .CLK(clk_bF$buf110),
    .D(_1521_[8]),
    .Q(\datapath_1.regfile_1.regOut[24] [8]),
    .R(rst_bF$buf58),
    .S(vdd)
);

AND2X2 _11108_ (
    .A(_1370_),
    .B(_1369_),
    .Y(_1323_[23])
);

FILL FILL_1__13611_ (
);

AND2X2 _15781_ (
    .A(_4135__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_4731_)
);

FILL FILL_0__15496_ (
);

FILL FILL401280x113620 (
);

OR2X2 _15361_ (
    .A(_4313_),
    .B(_4316_),
    .Y(_4317_)
);

FILL FILL452200x291460 (
);

FILL FILL_0__13809_ (
);

AND2X2 _16986_ (
    .A(_4151__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_5917_)
);

OR2X2 _16566_ (
    .A(_5500_),
    .B(_5503_),
    .Y(_5504_)
);

AND2X2 _16146_ (
    .A(_4183__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_5090_)
);

DFFSR _11281_ (
    .CLK(clk_bF$buf99),
    .D(_1389_[19]),
    .Q(\datapath_1.regfile_1.regOut[22] [19]),
    .R(rst_bF$buf19),
    .S(vdd)
);

FILL FILL_1__9418_ (
);

FILL FILL229520x286520 (
);

FILL FILL_0__17642_ (
);

OR2X2 _8488_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .B(_68__bF$buf3),
    .Y(_24_)
);

FILL FILL_1__10736_ (
);

FILL FILL352640x370500 (
);

INVX1 _12486_ (
    .A(\control_1.reg_state.dout [0]),
    .Y(_2091_)
);

DFFSR _12066_ (
    .CLK(clk_bF$buf7),
    .D(_1785_[30]),
    .Q(\datapath_1.regfile_1.regOut[28] [30]),
    .R(rst_bF$buf75),
    .S(vdd)
);

AND2X2 _18712_ (
    .A(_6302__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_7617_)
);

FILL FILL_0__18427_ (
);

FILL FILL_0__18007_ (
);

FILL FILL_0__13562_ (
);

FILL FILL_0__13142_ (
);

FILL FILL_0__8528_ (
);

FILL FILL61560x271700 (
);

FILL FILL453720x54340 (
);

AND2X2 _14632_ (
    .A(_3807_),
    .B(_3806_),
    .Y(_3804_[1])
);

OR2X2 _14212_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[23]),
    .Y(_3586_)
);

FILL FILL411160x88920 (
);

FILL FILL295640x187720 (
);

FILL FILL_0__18180_ (
);

FILL FILL433200x103740 (
);

FILL FILL_1__16559_ (
);

AND2X2 _15837_ (
    .A(_4217__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_4786_)
);

OR2X2 _15417_ (
    .A(_4341_),
    .B(_4372_),
    .Y(_4373_)
);

OR2X2 _10972_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .B(_1322__bF$buf0),
    .Y(_1300_)
);

FILL FILL_0__10687_ (
);

FILL FILL72200x143260 (
);

FILL FILL_0__10267_ (
);

FILL FILL_1__17500_ (
);

OR2X2 _10552_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .B(_1124__bF$buf3),
    .Y(_1080_)
);

DFFSR _10132_ (
    .CLK(clk_bF$buf57),
    .D(_795_[31]),
    .Q(\datapath_1.regfile_1.regOut[13] [31]),
    .R(rst_bF$buf81),
    .S(vdd)
);

FILL FILL_0__19385_ (
);

OR2X2 _19250_ (
    .A(_8143_),
    .B(_8146_),
    .Y(_8147_)
);

FILL FILL_1__12899_ (
);

DFFSR _8700_ (
    .CLK(clk_bF$buf3),
    .D(_69_[18]),
    .Q(\datapath_1.regfile_1.regOut[2] [18]),
    .R(rst_bF$buf58),
    .S(vdd)
);

FILL FILL_1__18705_ (
);

OR2X2 _11757_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_1703_)
);

FILL FILL51680x74100 (
);

OR2X2 _11337_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_1483_)
);

FILL FILL_0__12833_ (
);

FILL FILL259160x123500 (
);

FILL FILL384560x39520 (
);

OR2X2 _15590_ (
    .A(_4541_),
    .B(_4542_),
    .Y(_4543_)
);

AND2X2 _15170_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_4128_)
);

FILL FILL201400x281580 (
);

AND2X2 _9905_ (
    .A(_748_),
    .B(_747_),
    .Y(_729_[9])
);

FILL FILL445360x138320 (
);

FILL FILL432440x4940 (
);

FILL FILL_0__13618_ (
);

OR2X2 _13903_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.PCJump [29]),
    .Y(_3335_)
);

AND2X2 _16795_ (
    .A(_4200__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_5729_)
);

FILL FILL95760x24700 (
);

OR2X2 _16375_ (
    .A(_5315_),
    .B(_5308_),
    .Y(_5316_)
);

AND2X2 _11090_ (
    .A(_1358_),
    .B(_1357_),
    .Y(_1323_[17])
);

FILL FILL_0__17451_ (
);

FILL FILL_0__17031_ (
);

FILL FILL293360x370500 (
);

FILL FILL371640x93860 (
);

FILL FILL_1__10545_ (
);

BUFX2 BUFX2_insert590 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf49)
);

BUFX2 BUFX2_insert591 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf48)
);

BUFX2 BUFX2_insert592 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf47)
);

BUFX2 BUFX2_insert593 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf46)
);

BUFX2 BUFX2_insert594 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf45)
);

BUFX2 BUFX2_insert595 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf44)
);

BUFX2 BUFX2_insert596 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf43)
);

BUFX2 BUFX2_insert597 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf42)
);

BUFX2 BUFX2_insert598 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf41)
);

BUFX2 BUFX2_insert599 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf40)
);

DFFSR _12295_ (
    .CLK(clk_bF$buf63),
    .D(_1917_[1]),
    .Q(\datapath_1.regfile_1.regOut[30] [1]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL_0__18656_ (
);

OR2X2 _18941_ (
    .A(_7842_),
    .B(_7841_),
    .Y(_7843_)
);

OR2X2 _18521_ (
    .A(_7428_),
    .B(_7427_),
    .Y(_7429_)
);

FILL FILL281200x158080 (
);

OR2X2 _18101_ (
    .A(_7014_),
    .B(_7015_),
    .Y(_7016_)
);

FILL FILL_0__13791_ (
);

FILL FILL_0__13371_ (
);

OR2X2 _10608_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_1117_)
);

FILL FILL56240x4940 (
);

FILL FILL_1__15163_ (
);

FILL FILL206720x19760 (
);

OR2X2 _19306_ (
    .A(_8200_),
    .B(_8201_),
    .Y(_8202_)
);

FILL FILL300960x187720 (
);

DFFSR _14861_ (
    .CLK(clk_bF$buf58),
    .D(_3870_[9]),
    .Q(_2_[9]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__14576_ (
);

FILL FILL_0__14156_ (
);

OR2X2 _14441_ (
    .A(vdd),
    .B(\datapath_1.Data [24]),
    .Y(_3720_)
);

OR2X2 _14021_ (
    .A(_3437_),
    .B(_3436_),
    .Y(_3438_)
);

FILL FILL236360x266760 (
);

FILL FILL126920x34580 (
);

AND2X2 _15646_ (
    .A(_4195__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_4598_)
);

AND2X2 _15226_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_4184_)
);

AND2X2 _10781_ (
    .A(_1192_),
    .B(_1255_),
    .Y(_1191_[0])
);

FILL FILL_0__10076_ (
);

DFFSR _10361_ (
    .CLK(clk_bF$buf17),
    .D(_927_[2]),
    .Q(\datapath_1.regfile_1.regOut[15] [2]),
    .R(rst_bF$buf49),
    .S(vdd)
);

FILL FILL91200x123500 (
);

FILL FILL_0__16722_ (
);

FILL FILL_0__16302_ (
);

FILL FILL505400x59280 (
);

FILL FILL_0__9295_ (
);

OR2X2 _11986_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .B(_1850__bF$buf3),
    .Y(_1816_)
);

OR2X2 _11566_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .B(_1652__bF$buf3),
    .Y(_1596_)
);

DFFSR _11146_ (
    .CLK(clk_bF$buf106),
    .D(_1323_[13]),
    .Q(\datapath_1.regfile_1.regOut[21] [13]),
    .R(rst_bF$buf0),
    .S(vdd)
);

FILL FILL_0__17927_ (
);

FILL FILL_0__17507_ (
);

FILL FILL_0__12642_ (
);

FILL FILL133000x256880 (
);

FILL FILL316920x316160 (
);

DFFSR _9714_ (
    .CLK(clk_bF$buf60),
    .D(_597_[0]),
    .Q(\datapath_1.regfile_1.regOut[10] [0]),
    .R(rst_bF$buf101),
    .S(vdd)
);

FILL FILL156560x242060 (
);

FILL FILL494760x350740 (
);

FILL FILL_1__14014_ (
);

OR2X2 _13712_ (
    .A(_3188_),
    .B(_3189_),
    .Y(_3190_)
);

FILL FILL_0__13007_ (
);

FILL FILL234840x222300 (
);

OR2X2 _16184_ (
    .A(_5112_),
    .B(_5127_),
    .Y(_5128_)
);

FILL FILL173280x158080 (
);

FILL FILL_0__17680_ (
);

FILL FILL_1__15639_ (
);

FILL FILL_1__10354_ (
);

FILL FILL161880x34580 (
);

AND2X2 _14917_ (
    .A(_3957_),
    .B(_3956_),
    .Y(_3936_[10])
);

AND2X2 _17389_ (
    .A(_6296_),
    .B(_6204_),
    .Y(_6315_)
);

FILL FILL_1__19472_ (
);

FILL FILL74480x242060 (
);

AND2X2 _18750_ (
    .A(_6315__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [21]),
    .Y(_7655_)
);

FILL FILL_0__18465_ (
);

AND2X2 _18330_ (
    .A(_6326__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_7241_)
);

FILL FILL_0__18045_ (
);

FILL FILL378480x153140 (
);

FILL FILL_0__8986_ (
);

OR2X2 _10837_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .B(_1256__bF$buf1),
    .Y(_1230_)
);

OR2X2 _10417_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .B(_1058__bF$buf3),
    .Y(_1010_)
);

FILL FILL283480x113620 (
);

DFFSR _19535_ (
    .CLK(clk_bF$buf28),
    .D(_8320_[12]),
    .Q(\datapath_1.regfile_1.regOut[0] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

OR2X2 _19115_ (
    .A(_8006_),
    .B(_8013_),
    .Y(_8014_)
);

FILL FILL294880x182780 (
);

OR2X2 _14670_ (
    .A(\datapath_1.rd1 [14]),
    .B(_3869__bF$buf1),
    .Y(_3833_)
);

FILL FILL_0__14385_ (
);

OR2X2 _14250_ (
    .A(\datapath_1.ALUResult [3]),
    .B(_3671__bF$buf0),
    .Y(_3613_)
);

FILL FILL38000x9880 (
);

FILL FILL450680x286520 (
);

FILL FILL194560x276640 (
);

FILL FILL367840x296400 (
);

FILL FILL418000x207480 (
);

FILL FILL505400x212420 (
);

AND2X2 _15875_ (
    .A(_4208__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_4823_)
);

OR2X2 _15455_ (
    .A(_4408_),
    .B(_4409_),
    .Y(_4410_)
);

INVX1 _15035_ (
    .A(_4023_),
    .Y(_4024_)
);

OR2X2 _10590_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_1105_)
);

OR2X2 _10170_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_885_)
);

FILL FILL_0__16951_ (
);

FILL FILL_0__16531_ (
);

FILL FILL_0__16111_ (
);

FILL FILL448400x163020 (
);

DFFSR _11795_ (
    .CLK(clk_bF$buf11),
    .D(_1653_[17]),
    .Q(\datapath_1.regfile_1.regOut[26] [17]),
    .R(rst_bF$buf36),
    .S(vdd)
);

FILL FILL_1__18323_ (
);

AND2X2 _11375_ (
    .A(_1508_),
    .B(_1507_),
    .Y(_1455_[26])
);

FILL FILL60800x281580 (
);

FILL FILL257640x316160 (
);

OR2X2 _17601_ (
    .A(_6516_),
    .B(_6523_),
    .Y(_6524_)
);

FILL FILL_0__12871_ (
);

FILL FILL364800x192660 (
);

OR2X2 _9943_ (
    .A(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .B(_794__bF$buf1),
    .Y(_774_)
);

OR2X2 _9523_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .B(_596__bF$buf1),
    .Y(_554_)
);

OR2X2 _9103_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(_398__bF$buf4),
    .Y(_334_)
);

FILL FILL_1__14663_ (
);

AND2X2 _18806_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_7710_)
);

FILL FILL_0_BUFX2_insert230 (
);

FILL FILL_0_BUFX2_insert231 (
);

FILL FILL_0_BUFX2_insert232 (
);

FILL FILL_0_BUFX2_insert233 (
);

FILL FILL367080x311220 (
);

OR2X2 _13941_ (
    .A(_3367_),
    .B(_3368_),
    .Y(_3369_)
);

FILL FILL_0__13656_ (
);

FILL FILL_0__13236_ (
);

FILL FILL_0_BUFX2_insert235 (
);

AND2X2 _13521_ (
    .A(_3035_),
    .B(_3034_),
    .Y(_1_[10])
);

NAND2X1 _13101_ (
    .A(_2524_),
    .B(_2654_),
    .Y(_2655_)
);

FILL FILL_0_BUFX2_insert237 (
);

FILL FILL_0_BUFX2_insert239 (
);

FILL FILL38760x256880 (
);

FILL FILL_1__9265_ (
);

BUFX2 BUFX2_insert1150 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf4 )
);

BUFX2 BUFX2_insert1151 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf3 )
);

BUFX2 BUFX2_insert1152 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf2 )
);

BUFX2 BUFX2_insert1153 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf1 )
);

BUFX2 BUFX2_insert1154 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf0 )
);

BUFX2 BUFX2_insert1155 (
    .A(_3347_),
    .Y(_3347__bF$buf4)
);

BUFX2 BUFX2_insert1156 (
    .A(_3347_),
    .Y(_3347__bF$buf3)
);

BUFX2 BUFX2_insert1157 (
    .A(_3347_),
    .Y(_3347__bF$buf2)
);

BUFX2 BUFX2_insert1158 (
    .A(_3347_),
    .Y(_3347__bF$buf1)
);

FILL FILL_1__15028_ (
);

BUFX2 BUFX2_insert1159 (
    .A(_3347_),
    .Y(_3347__bF$buf0)
);

FILL FILL444600x44460 (
);

FILL FILL_1__10163_ (
);

DFFSR _14726_ (
    .CLK(clk_bF$buf4),
    .D(_3804_[3]),
    .Q(\datapath_1.a [3]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _14306_ (
    .A(vdd),
    .B(ALUOut[22]),
    .Y(_3650_)
);

FILL FILL410400x316160 (
);

BUFX2 BUFX2_insert970 (
    .A(_4197_),
    .Y(_4197__bF$buf0)
);

BUFX2 BUFX2_insert971 (
    .A(_1190_),
    .Y(_1190__bF$buf4)
);

BUFX2 BUFX2_insert972 (
    .A(_1190_),
    .Y(_1190__bF$buf3)
);

BUFX2 BUFX2_insert973 (
    .A(_1190_),
    .Y(_1190__bF$buf2)
);

FILL FILL20520x54340 (
);

BUFX2 BUFX2_insert974 (
    .A(_1190_),
    .Y(_1190__bF$buf1)
);

BUFX2 BUFX2_insert975 (
    .A(_1190_),
    .Y(_1190__bF$buf0)
);

BUFX2 BUFX2_insert976 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf4 )
);

OR2X2 _17198_ (
    .A(_6124_),
    .B(_6125_),
    .Y(_6126_)
);

BUFX2 BUFX2_insert977 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf3 )
);

FILL FILL_0__15802_ (
);

BUFX2 BUFX2_insert978 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf2 )
);

BUFX2 BUFX2_insert979 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf1 )
);

FILL FILL127680x64220 (
);

FILL FILL_0__18274_ (
);

FILL FILL414200x237120 (
);

FILL FILL205960x123500 (
);

DFFSR _10646_ (
    .CLK(clk_bF$buf53),
    .D(_1059_[29]),
    .Q(\datapath_1.regfile_1.regOut[17] [29]),
    .R(rst_bF$buf6),
    .S(vdd)
);

AND2X2 _10226_ (
    .A(_922_),
    .B(_921_),
    .Y(_861_[30])
);

FILL FILL_0__11302_ (
);

FILL FILL_0__19479_ (
);

OR2X2 _19344_ (
    .A(_8238_),
    .B(_8239_),
    .Y(_8240_)
);

FILL FILL_0__14194_ (
);

FILL FILL281200x311220 (
);

FILL FILL183920x69160 (
);

FILL FILL503880x98800 (
);

FILL FILL72200x306280 (
);

FILL FILL_0__12927_ (
);

FILL FILL_0__12507_ (
);

FILL FILL376200x217360 (
);

OR2X2 _15684_ (
    .A(_4633_),
    .B(_4634_),
    .Y(_4635_)
);

AND2X2 _15264_ (
    .A(_4127_),
    .B(_4171_),
    .Y(_4222_)
);

FILL FILL82840x0 (
);

FILL FILL_0__16760_ (
);

FILL FILL17480x276640 (
);

FILL FILL62320x251940 (
);

FILL FILL53960x128440 (
);

FILL FILL148960x88920 (
);

OR2X2 _16889_ (
    .A(_5821_),
    .B(_5790_),
    .Y(_5822_)
);

AND2X2 _16469_ (
    .A(_4197__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_5408_)
);

AND2X2 _16049_ (
    .A(_4189__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_4995_)
);

FILL FILL_1__18972_ (
);

OR2X2 _11184_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_1401_)
);

FILL FILL357960x360620 (
);

FILL FILL_0__17545_ (
);

OR2X2 _17830_ (
    .A(_6748_),
    .B(_6735_),
    .Y(_6749_)
);

AND2X2 _17410_ (
    .A(_6335_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd1 [0])
);

FILL FILL_0__17125_ (
);

FILL FILL_0__12680_ (
);

FILL FILL458280x247000 (
);

FILL FILL488680x158080 (
);

AND2X2 _9752_ (
    .A(_666_),
    .B(_665_),
    .Y(_663_[1])
);

DFFSR _9332_ (
    .CLK(clk_bF$buf36),
    .D(_399_[5]),
    .Q(\datapath_1.regfile_1.regOut[7] [5]),
    .R(rst_bF$buf25),
    .S(vdd)
);

AND2X2 _12389_ (
    .A(_2024_),
    .B(_2023_),
    .Y(_1983_[20])
);

FILL FILL_1__14052_ (
);

FILL FILL374680x276640 (
);

AND2X2 _18615_ (
    .A(_6255__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_7522_)
);

FILL FILL_0__13885_ (
);

OR2X2 _13750_ (
    .A(_3222_),
    .B(_3221_),
    .Y(_3223_)
);

NAND2X1 _13330_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2871_)
);

FILL FILL133760x311220 (
);

FILL FILL368600x232180 (
);

FILL FILL299440x44460 (
);

FILL FILL483360x44460 (
);

FILL FILL_1__15677_ (
);

OR2X2 _14955_ (
    .A(\datapath_1.mux_pcsrc.dout [23]),
    .B(_4001__bF$buf1),
    .Y(_3983_)
);

OR2X2 _14535_ (
    .A(memoryOutData[12]),
    .B(_3803__bF$buf0),
    .Y(_3763_)
);

AND2X2 _14115_ (
    .A(_3347__bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3518_)
);

FILL FILL254600x350740 (
);

FILL FILL_0__15611_ (
);

FILL FILL_0__18083_ (
);

FILL FILL_1__11597_ (
);

FILL FILL258400x271700 (
);

FILL FILL51680x311220 (
);

DFFSR _10875_ (
    .CLK(clk_bF$buf41),
    .D(_1191_[0]),
    .Q(\datapath_1.regfile_1.regOut[19] [0]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL_1__17823_ (
);

OR2X2 _10455_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_1035_)
);

OR2X2 _10035_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_815_)
);

FILL FILL_0__16816_ (
);

OR2X2 _19153_ (
    .A(_8048_),
    .B(_8051_),
    .Y(_8052_)
);

AND2X2 _8603_ (
    .A(_80_),
    .B(_79_),
    .Y(_69_[5])
);

FILL FILL285760x227240 (
);

FILL FILL495520x103740 (
);

FILL FILL_0__9389_ (
);

FILL FILL164160x4940 (
);

FILL FILL_0__12736_ (
);

FILL FILL234080x74100 (
);

NAND2X1 _12601_ (
    .A(_2163_),
    .B(_2165_),
    .Y(_2166_)
);

FILL FILL166440x49400 (
);

FILL FILL212040x118560 (
);

AND2X2 _15493_ (
    .A(_4160__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_4447_)
);

NAND2X1 _15073_ (
    .A(_4024_),
    .B(_4059_),
    .Y(_4060_)
);

OR2X2 _9808_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .B(_728__bF$buf1),
    .Y(_704_)
);

FILL FILL430160x242060 (
);

FILL FILL320720x330980 (
);

OR2X2 _13806_ (
    .A(_3270_),
    .B(_3269_),
    .Y(_3271_)
);

FILL FILL408120x222300 (
);

AND2X2 _16698_ (
    .A(_5633_),
    .B(_4065__bF$buf5),
    .Y(\datapath_1.rd2 [22])
);

OR2X2 _16278_ (
    .A(_5219_),
    .B(_5218_),
    .Y(_5220_)
);

FILL FILL129960x113620 (
);

FILL FILL_0__17774_ (
);

FILL FILL263720x281580 (
);

FILL FILL_1__10448_ (
);

DFFSR _9981_ (
    .CLK(clk_bF$buf24),
    .D(_729_[9]),
    .Q(\datapath_1.regfile_1.regOut[12] [9]),
    .R(rst_bF$buf83),
    .S(vdd)
);

OR2X2 _9561_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_579_)
);

OR2X2 _9141_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_359_)
);

FILL FILL224200x345800 (
);

INVX2 _12198_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .Y(_1982_)
);

FILL FILL_1__19146_ (
);

FILL FILL_0__18979_ (
);

AND2X2 _18844_ (
    .A(_6271__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_7747_)
);

FILL FILL_0_BUFX2_insert610 (
);

FILL FILL260680x326040 (
);

FILL FILL_0_BUFX2_insert611 (
);

FILL FILL_0__18139_ (
);

AND2X2 _18424_ (
    .A(_6259__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_7334_)
);

FILL FILL297920x64220 (
);

FILL FILL_0_BUFX2_insert612 (
);

AND2X2 _18004_ (
    .A(_6317__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_6920_)
);

FILL FILL_0_BUFX2_insert613 (
);

FILL FILL_0__13274_ (
);

FILL FILL_0_BUFX2_insert615 (
);

FILL FILL470440x202540 (
);

FILL FILL_0_BUFX2_insert617 (
);

FILL FILL_0_BUFX2_insert619 (
);

FILL FILL64600x138320 (
);

OR2X2 _19209_ (
    .A(_8103_),
    .B(_8106_),
    .Y(_8107_)
);

AND2X2 _14764_ (
    .A(_3875_),
    .B(_3874_),
    .Y(_3870_[2])
);

FILL FILL_0__14059_ (
);

DFFSR _14344_ (
    .CLK(clk_bF$buf50),
    .D(_3606_[8]),
    .Q(ALUOut[8]),
    .R(rst_bF$buf18),
    .S(vdd)
);

FILL FILL_0__15420_ (
);

FILL FILL385320x286520 (
);

AND2X2 _15969_ (
    .A(_4200__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_4916_)
);

OR2X2 _15549_ (
    .A(_4500_),
    .B(_4501_),
    .Y(_4502_)
);

AND2X2 _15129_ (
    .A(_4100_),
    .B(_4104_),
    .Y(_4105_)
);

OR2X2 _10684_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .B(_1190__bF$buf2),
    .Y(_1148_)
);

FILL FILL_0__10399_ (
);

OR2X2 _10264_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(_992__bF$buf2),
    .Y(_928_)
);

FILL FILL_0__16625_ (
);

AND2X2 _16910_ (
    .A(_4135__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_5842_)
);

FILL FILL_0__11760_ (
);

FILL FILL_0__11340_ (
);

AND2X2 _19382_ (
    .A(_6229__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_8277_)
);

FILL FILL_0__19097_ (
);

DFFSR _8832_ (
    .CLK(clk_bF$buf1),
    .D(_135_[21]),
    .Q(\datapath_1.regfile_1.regOut[3] [21]),
    .R(rst_bF$buf38),
    .S(vdd)
);

BUFX2 _8412_ (
    .A(_1_[20]),
    .Y(memoryAddress[20])
);

FILL FILL_1__18837_ (
);

OR2X2 _11889_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_1771_)
);

OR2X2 _11469_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_1551_)
);

OR2X2 _11049_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_1331_)
);

FILL FILL_1__13552_ (
);

FILL FILL_1__13132_ (
);

OR2X2 _12830_ (
    .A(_2394_),
    .B(_2391_),
    .Y(_2395_)
);

FILL FILL_0__12125_ (
);

AND2X2 _12410_ (
    .A(_2038_),
    .B(_2037_),
    .Y(_1983_[27])
);

FILL FILL155800x256880 (
);

OR2X2 _9617_ (
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .Y(_661_)
);

AND2X2 _13615_ (
    .A(_3087__bF$buf2),
    .B(\datapath_1.ALUResult [3]),
    .Y(_3107_)
);

OR2X2 _16087_ (
    .A(_5031_),
    .B(_5028_),
    .Y(_5032_)
);

FILL FILL_1__9359_ (
);

FILL FILL113240x158080 (
);

FILL FILL_0__17583_ (
);

FILL FILL_0__17163_ (
);

FILL FILL168720x4940 (
);

OR2X2 _9790_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .B(_728__bF$buf4),
    .Y(_692_)
);

OR2X2 _9370_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .B(_530__bF$buf3),
    .Y(_472_)
);

FILL FILL79040x330980 (
);

FILL FILL_0__10611_ (
);

FILL FILL_0__18788_ (
);

AND2X2 _18653_ (
    .A(_6250__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_7559_)
);

FILL FILL_0__18368_ (
);

FILL FILL118560x54340 (
);

OR2X2 _18233_ (
    .A(_7145_),
    .B(_7144_),
    .Y(_7146_)
);

FILL FILL_0__13083_ (
);

FILL FILL234840x29640 (
);

FILL FILL_0__8469_ (
);

FILL FILL248520x158080 (
);

FILL FILL409640x39520 (
);

FILL FILL309320x128440 (
);

FILL FILL_0__9830_ (
);

FILL FILL_0__11816_ (
);

FILL FILL_0__9410_ (
);

FILL FILL31160x158080 (
);

AND2X2 _19438_ (
    .A(_8327_),
    .B(_8326_),
    .Y(_8320_[3])
);

AND2X2 _19018_ (
    .A(_6312__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_7919_)
);

DFFSR _14993_ (
    .CLK(clk_bF$buf20),
    .D(_3936_[12]),
    .Q(\datapath_1.mux_iord.din0 [12]),
    .R(rst_bF$buf29),
    .S(vdd)
);

OR2X2 _14573_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_3788_)
);

OR2X2 _14153_ (
    .A(\datapath_1.Data [3]),
    .B(_3605__bF$buf2),
    .Y(_3547_)
);

FILL FILL151240x59280 (
);

AND2X2 _15778_ (
    .A(_4241__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_4728_)
);

AND2X2 _15358_ (
    .A(_4151__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_4314_)
);

FILL FILL_1__17441_ (
);

DFFSR _10493_ (
    .CLK(clk_bF$buf29),
    .D(_993_[5]),
    .Q(\datapath_1.regfile_1.regOut[16] [5]),
    .R(rst_bF$buf40),
    .S(vdd)
);

AND2X2 _10073_ (
    .A(_840_),
    .B(_839_),
    .Y(_795_[22])
);

FILL FILL358720x113620 (
);

FILL FILL_0__16014_ (
);

OR2X2 _19191_ (
    .A(_8088_),
    .B(_8087_),
    .Y(_8089_)
);

FILL FILL288800x118560 (
);

OR2X2 _8641_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .B(_134__bF$buf1),
    .Y(_106_)
);

OR2X2 _11698_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .B(_1718__bF$buf4),
    .Y(_1664_)
);

DFFSR _11278_ (
    .CLK(clk_bF$buf53),
    .D(_1389_[16]),
    .Q(\datapath_1.regfile_1.regOut[22] [16]),
    .R(rst_bF$buf73),
    .S(vdd)
);

FILL FILL_1__13781_ (
);

OR2X2 _17924_ (
    .A(_6841_),
    .B(_6840_),
    .Y(_6842_)
);

FILL FILL_0__17639_ (
);

FILL FILL_0__17219_ (
);

OR2X2 _17504_ (
    .A(_6420_),
    .B(_6427_),
    .Y(_6428_)
);

FILL FILL_0__12774_ (
);

DFFSR _9846_ (
    .CLK(clk_bF$buf44),
    .D(_663_[3]),
    .Q(\datapath_1.regfile_1.regOut[11] [3]),
    .R(rst_bF$buf97),
    .S(vdd)
);

OR2X2 _9426_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_509_)
);

OR2X2 _9006_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_289_)
);

FILL FILL66880x237120 (
);

FILL FILL389880x311220 (
);

OR2X2 _18709_ (
    .A(_7581_),
    .B(_7614_),
    .Y(_7615_)
);

FILL FILL56240x197600 (
);

FILL FILL_0__13979_ (
);

OR2X2 _13844_ (
    .A(\datapath_1.a [9]),
    .B(_3342__bF$buf3),
    .Y(_3296_)
);

FILL FILL_0__13139_ (
);

NOR2X1 _13424_ (
    .A(_2854_),
    .B(_2852_),
    .Y(_2959_)
);

NOR2X1 _13004_ (
    .A(_2501_),
    .B(_2318_),
    .Y(_2564_)
);

FILL FILL_0__14500_ (
);

FILL FILL237120x316160 (
);

FILL FILL_1__9168_ (
);

FILL FILL324520x321100 (
);

FILL FILL_0__17392_ (
);

FILL FILL_1__10486_ (
);

AND2X2 _14629_ (
    .A(_3805_),
    .B(_3868_),
    .Y(_3804_[0])
);

OR2X2 _14209_ (
    .A(MemToReg_bF$buf0),
    .B(ALUOut[22]),
    .Y(_3584_)
);

FILL FILL410400x54340 (
);

FILL FILL_0__10840_ (
);

FILL FILL_0__10420_ (
);

AND2X2 _18882_ (
    .A(_6236__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_7785_)
);

FILL FILL_0__18597_ (
);

AND2X2 _18462_ (
    .A(_6317__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_7371_)
);

FILL FILL431680x93860 (
);

NOR2X1 _18042_ (
    .A(_6310__bF$buf4),
    .B(_6957_),
    .Y(_6958_)
);

FILL FILL350360x128440 (
);

OR2X2 _10969_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .B(_1322__bF$buf2),
    .Y(_1298_)
);

FILL FILL_1__17917_ (
);

OR2X2 _10549_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_1124__bF$buf3),
    .Y(_1078_)
);

DFFSR _10129_ (
    .CLK(clk_bF$buf74),
    .D(_795_[28]),
    .Q(\datapath_1.regfile_1.regOut[13] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _11910_ (
    .CLK(clk_bF$buf44),
    .D(_1719_[3]),
    .Q(\datapath_1.regfile_1.regOut[27] [3]),
    .R(rst_bF$buf16),
    .S(vdd)
);

FILL FILL_0__11625_ (
);

FILL FILL_0__11205_ (
);

AND2X2 _19247_ (
    .A(_6264__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_8144_)
);

FILL FILL373160x212420 (
);

FILL FILL478040x34580 (
);

FILL FILL_0__14097_ (
);

OR2X2 _14382_ (
    .A(memoryOutData[4]),
    .B(_3737__bF$buf3),
    .Y(_3681_)
);

FILL FILL_1__13417_ (
);

FILL FILL345040x345800 (
);

OR2X2 _15587_ (
    .A(_4538_),
    .B(_4539_),
    .Y(_4540_)
);

NOR2X1 _15167_ (
    .A(_4124_),
    .B(_4065__bF$buf6),
    .Y(\datapath_1.regfile_1.regEn [31])
);

FILL FILL_1__8859_ (
);

FILL FILL_0__16663_ (
);

FILL FILL_0__16243_ (
);

AND2X2 _8870_ (
    .A(_218_),
    .B(_217_),
    .Y(_201_[8])
);

BUFX2 _8450_ (
    .A(_2_[26]),
    .Y(memoryWriteData[26])
);

AND2X2 _11087_ (
    .A(_1356_),
    .B(_1355_),
    .Y(_1323_[16])
);

FILL FILL_1__13170_ (
);

FILL FILL_0__17868_ (
);

FILL FILL_0__17448_ (
);

OR2X2 _17733_ (
    .A(_6622_),
    .B(_6653_),
    .Y(_6654_)
);

FILL FILL88920x172900 (
);

AND2X2 _17313_ (
    .A(_6238__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_6239_)
);

FILL FILL403560x113620 (
);

FILL FILL_0__12583_ (
);

FILL FILL414960x182780 (
);

OR2X2 _9655_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .B(_662__bF$buf0),
    .Y(_622_)
);

OR2X2 _9235_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .B(_464__bF$buf1),
    .Y(_402_)
);

FILL FILL10640x365560 (
);

FILL FILL_0__8910_ (
);

FILL FILL_1__14795_ (
);

OR2X2 _18938_ (
    .A(_7838_),
    .B(_7839_),
    .Y(_7840_)
);

OR2X2 _18518_ (
    .A(_7425_),
    .B(_7424_),
    .Y(_7426_)
);

FILL FILL295640x232180 (
);

FILL FILL_0__13788_ (
);

FILL FILL_0__13368_ (
);

OR2X2 _13653_ (
    .A(_3139_),
    .B(_3136_),
    .Y(\datapath_1.mux_pcsrc.dout [8])
);

XOR2X1 _13233_ (
    .A(_2215_),
    .B(_2730_),
    .Y(_2779_)
);

FILL FILL288800x54340 (
);

FILL FILL_1__10295_ (
);

DFFSR _14858_ (
    .CLK(clk_bF$buf77),
    .D(_3870_[6]),
    .Q(_2_[6]),
    .R(rst_bF$buf65),
    .S(vdd)
);

OR2X2 _14438_ (
    .A(vdd),
    .B(\datapath_1.Data [23]),
    .Y(_3718_)
);

FILL FILL354920x370500 (
);

OR2X2 _14018_ (
    .A(_3433_),
    .B(_3434_),
    .Y(_3435_)
);

FILL FILL65360x103740 (
);

FILL FILL_1__16941_ (
);

FILL FILL_1__16521_ (
);

FILL FILL_0_CLKBUF1_insert220 (
);

FILL FILL_0_CLKBUF1_insert221 (
);

FILL FILL300200x103740 (
);

FILL FILL_0__15514_ (
);

FILL FILL_0_CLKBUF1_insert223 (
);

OR2X2 _18691_ (
    .A(_7589_),
    .B(_7596_),
    .Y(_7597_)
);

AND2X2 _18271_ (
    .A(_6216__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_7183_)
);

FILL FILL63840x271700 (
);

OR2X2 _10778_ (
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .Y(_1255_)
);

AND2X2 _10358_ (
    .A(_990_),
    .B(_989_),
    .Y(_927_[31])
);

FILL FILL_1__17306_ (
);

FILL FILL_0__11434_ (
);

OR2X2 _19476_ (
    .A(gnd),
    .B(_8385__bF$buf0),
    .Y(_8353_)
);

OR2X2 _19056_ (
    .A(_7952_),
    .B(_7955_),
    .Y(_7956_)
);

OR2X2 _14191_ (
    .A(MemToReg_bF$buf3),
    .B(ALUOut[16]),
    .Y(_3572_)
);

FILL FILL2280x187720 (
);

OR2X2 _8926_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .B(_266__bF$buf3),
    .Y(_256_)
);

FILL FILL297920x187720 (
);

OR2X2 _8506_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .B(_68__bF$buf3),
    .Y(_36_)
);

FILL FILL_1__13646_ (
);

FILL FILL_1_BUFX2_insert541 (
);

AND2X2 _12924_ (
    .A(_2486_),
    .B(_2488_),
    .Y(_2489_)
);

FILL FILL_0__12639_ (
);

FILL FILL_1_BUFX2_insert543 (
);

FILL FILL_0__12219_ (
);

NAND2X1 _12504_ (
    .A(\control_1.reg_state.dout [2]),
    .B(_2100_),
    .Y(_2101_)
);

FILL FILL_1_BUFX2_insert545 (
);

AND2X2 _15396_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_4352_)
);

FILL FILL_0__16892_ (
);

FILL FILL_0__16472_ (
);

FILL FILL503120x172900 (
);

FILL FILL_0__16052_ (
);

FILL FILL40280x202540 (
);

OR2X2 _13709_ (
    .A(_3187_),
    .B(_3184_),
    .Y(\datapath_1.mux_pcsrc.dout [16])
);

FILL FILL19760x69160 (
);

FILL FILL_1__18264_ (
);

FILL FILL355680x182780 (
);

AND2X2 _17962_ (
    .A(_6271__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_6879_)
);

AND2X2 _17542_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_6465_)
);

FILL FILL_0__17257_ (
);

AND2X2 _17122_ (
    .A(_4172__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_6051_)
);

FILL FILL44080x123500 (
);

FILL FILL_0__12392_ (
);

FILL FILL447640x138320 (
);

AND2X2 _9884_ (
    .A(_734_),
    .B(_733_),
    .Y(_729_[2])
);

DFFSR _9464_ (
    .CLK(clk_bF$buf74),
    .D(_465_[8]),
    .Q(\datapath_1.regfile_1.regOut[8] [8]),
    .R(rst_bF$buf11),
    .S(vdd)
);

AND2X2 _9044_ (
    .A(_314_),
    .B(_313_),
    .Y(_267_[23])
);

FILL FILL_0__10705_ (
);

OR2X2 _18747_ (
    .A(_7651_),
    .B(_7650_),
    .Y(_7652_)
);

FILL FILL278160x360620 (
);

OR2X2 _18327_ (
    .A(_7235_),
    .B(_7237_),
    .Y(_7238_)
);

FILL FILL_0__13597_ (
);

OR2X2 _13882_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.mux_iord.din0 [22]),
    .Y(_3321_)
);

FILL FILL_0__13177_ (
);

AND2X2 _13462_ (
    .A(_2789_),
    .B(_2819_),
    .Y(_2995_)
);

INVX1 _13042_ (
    .A(_2599_),
    .Y(\datapath_1.ALUResult [24])
);

FILL FILL131480x133380 (
);

FILL FILL280440x24700 (
);

FILL FILL_0__19403_ (
);

FILL FILL464360x375440 (
);

FILL FILL295640x370500 (
);

FILL FILL_0__9924_ (
);

FILL FILL_0__9504_ (
);

FILL FILL204440x247000 (
);

OR2X2 _14667_ (
    .A(\datapath_1.rd1 [13]),
    .B(_3869__bF$buf1),
    .Y(_3831_)
);

OR2X2 _14247_ (
    .A(\datapath_1.ALUResult [2]),
    .B(_3671__bF$buf1),
    .Y(_3611_)
);

FILL FILL_0__15743_ (
);

FILL FILL53200x163020 (
);

FILL FILL95760x98800 (
);

OR2X2 _18080_ (
    .A(_6993_),
    .B(_6994_),
    .Y(_6995_)
);

FILL FILL504640x44460 (
);

OR2X2 _10587_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_1103_)
);

OR2X2 _10167_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_883_)
);

FILL FILL_1__12670_ (
);

FILL FILL_0__16528_ (
);

AND2X2 _16813_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_5747_)
);

FILL FILL_0__16108_ (
);

AND2X2 _19285_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_8182_)
);

FILL FILL207480x79040 (
);

AND2X2 _8735_ (
    .A(_148_),
    .B(_147_),
    .Y(_135_[6])
);

FILL FILL149720x34580 (
);

FILL FILL_0__12868_ (
);

OR2X2 _12733_ (
    .A(_2280_),
    .B(_2297_),
    .Y(_2298_)
);

DFFSR _12313_ (
    .CLK(clk_bF$buf19),
    .D(_1917_[19]),
    .Q(\datapath_1.regfile_1.regOut[30] [19]),
    .R(rst_bF$buf13),
    .S(vdd)
);

FILL FILL_0__12028_ (
);

FILL FILL126160x34580 (
);

FILL FILL34960x39520 (
);

FILL FILL435480x29640 (
);

OR2X2 _13938_ (
    .A(_3366_),
    .B(_3363_),
    .Y(\datapath_1.alu_1.ALUInB [2])
);

AND2X2 _13518_ (
    .A(_3033_),
    .B(_3032_),
    .Y(_1_[9])
);

FILL FILL_1__18493_ (
);

FILL FILL_0__17486_ (
);

AND2X2 _17771_ (
    .A(_6328__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_6691_)
);

FILL FILL_0__17066_ (
);

AND2X2 _17351_ (
    .A(_6275_),
    .B(_6276_),
    .Y(_6277_)
);

FILL FILL158840x242060 (
);

FILL FILL323000x148200 (
);

OR2X2 _9693_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_647_)
);

FILL FILL_1__16806_ (
);

FILL FILL232560x207480 (
);

OR2X2 _9273_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_427_)
);

FILL FILL_1__19278_ (
);

FILL FILL264480x19760 (
);

OR2X2 _18976_ (
    .A(_7875_),
    .B(_7876_),
    .Y(_7877_)
);

OR2X2 _18556_ (
    .A(_7462_),
    .B(_7463_),
    .Y(_7464_)
);

AND2X2 _18136_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_7050_)
);

OR2X2 _13691_ (
    .A(_3170_),
    .B(_3171_),
    .Y(_3172_)
);

AND2X2 _13271_ (
    .A(_2812_),
    .B(_2814_),
    .Y(_2815_)
);

FILL FILL38760x39520 (
);

FILL FILL175560x158080 (
);

FILL FILL_0__19212_ (
);

FILL FILL262960x163020 (
);

FILL FILL439280x29640 (
);

FILL FILL_0__11719_ (
);

FILL FILL_1__15198_ (
);

AND2X2 _14896_ (
    .A(_3943_),
    .B(_3942_),
    .Y(_3936_[3])
);

DFFSR _14476_ (
    .CLK(clk_bF$buf23),
    .D(_3672_[11]),
    .Q(\datapath_1.Data [11]),
    .R(rst_bF$buf22),
    .S(vdd)
);

OR2X2 _14056_ (
    .A(_3467_),
    .B(_3466_),
    .Y(_3468_)
);

FILL FILL76760x242060 (
);

FILL FILL_0__15132_ (
);

FILL FILL76000x340860 (
);

FILL FILL494000x227240 (
);

OR2X2 _10396_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .B(_1058__bF$buf3),
    .Y(_996_)
);

FILL FILL435480x276640 (
);

FILL FILL_0__16757_ (
);

OR2X2 _16622_ (
    .A(_5557_),
    .B(_5558_),
    .Y(_5559_)
);

FILL FILL_0__16337_ (
);

AND2X2 _16202_ (
    .A(_4234__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_5145_)
);

FILL FILL_0__11892_ (
);

FILL FILL_0__11472_ (
);

OR2X2 _19094_ (
    .A(_7993_),
    .B(_7992_),
    .Y(_7994_)
);

FILL FILL458280x360620 (
);

FILL FILL196840x276640 (
);

DFFSR _8964_ (
    .CLK(clk_bF$buf35),
    .D(_201_[24]),
    .Q(\datapath_1.regfile_1.regOut[4] [24]),
    .R(rst_bF$buf34),
    .S(vdd)
);

OR2X2 _8544_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_61_)
);

FILL FILL_1__18129_ (
);

OR2X2 _17827_ (
    .A(_6745_),
    .B(_6744_),
    .Y(_6746_)
);

OR2X2 _17407_ (
    .A(_6332_),
    .B(_6306_),
    .Y(_6333_)
);

FILL FILL_1_BUFX2_insert921 (
);

NAND3X1 _12962_ (
    .A(_2363_),
    .B(_2366_),
    .C(_2524_),
    .Y(_2525_)
);

FILL FILL_1_BUFX2_insert923 (
);

FILL FILL_0__12257_ (
);

AND2X2 _12542_ (
    .A(_2129_),
    .B(_2130_),
    .Y(_2131_)
);

AND2X2 _12122_ (
    .A(_1886_),
    .B(_1885_),
    .Y(_1851_[17])
);

FILL FILL_1_BUFX2_insert925 (
);

FILL FILL_0__18903_ (
);

AND2X2 _9749_ (
    .A(_664_),
    .B(_727_),
    .Y(_663_[0])
);

FILL FILL501600x365560 (
);

DFFSR _9329_ (
    .CLK(clk_bF$buf111),
    .D(_399_[2]),
    .Q(\datapath_1.regfile_1.regOut[7] [2]),
    .R(rst_bF$buf108),
    .S(vdd)
);

FILL FILL_0__16090_ (
);

FILL FILL226480x49400 (
);

FILL FILL319200x271700 (
);

OR2X2 _13747_ (
    .A(_3218_),
    .B(_3219_),
    .Y(_3220_)
);

INVX1 _13327_ (
    .A(_2410_),
    .Y(_2868_)
);

FILL FILL_1__15410_ (
);

FILL FILL416480x222300 (
);

FILL FILL505400x286520 (
);

FILL FILL_0__14823_ (
);

FILL FILL_0__14403_ (
);

FILL FILL486400x242060 (
);

NOR2X1 _17580_ (
    .A(_6310__bF$buf0),
    .B(_6502_),
    .Y(_6503_)
);

OR2X2 _17160_ (
    .A(_6087_),
    .B(_6084_),
    .Y(_6088_)
);

FILL FILL109440x88920 (
);

FILL FILL440040x44460 (
);

DFFSR _9082_ (
    .CLK(clk_bF$buf37),
    .D(_267_[13]),
    .Q(\datapath_1.regfile_1.regOut[5] [13]),
    .R(rst_bF$buf46),
    .S(vdd)
);

FILL FILL285000x355680 (
);

FILL FILL372400x360620 (
);

FILL FILL_1__11750_ (
);

FILL FILL_0__15608_ (
);

FILL FILL177080x128440 (
);

OR2X2 _18785_ (
    .A(_7687_),
    .B(_7688_),
    .Y(_7689_)
);

OR2X2 _18365_ (
    .A(_7275_),
    .B(_7272_),
    .Y(_7276_)
);

FILL FILL232560x345800 (
);

INVX1 _13080_ (
    .A(_2274_),
    .Y(_2635_)
);

FILL FILL_0__19021_ (
);

FILL FILL_1__12115_ (
);

FILL FILL_0__9962_ (
);

FILL FILL_0__11948_ (
);

FILL FILL_0__9542_ (
);

AND2X2 _11813_ (
    .A(_1720_),
    .B(_1783_),
    .Y(_1719_[0])
);

FILL FILL_0__11108_ (
);

FILL FILL313120x212420 (
);

OR2X2 _14285_ (
    .A(vdd),
    .B(ALUOut[15]),
    .Y(_3636_)
);

FILL FILL_0__15781_ (
);

FILL FILL324520x281580 (
);

FILL FILL_0__15361_ (
);

FILL FILL_0__16986_ (
);

FILL FILL_0__16566_ (
);

OR2X2 _16851_ (
    .A(_5782_),
    .B(_5783_),
    .Y(_5784_)
);

OR2X2 _16431_ (
    .A(_5370_),
    .B(_5367_),
    .Y(_5371_)
);

AND2X2 _16011_ (
    .A(_4160__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_4957_)
);

OR2X2 _8773_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .B(_200__bF$buf4),
    .Y(_174_)
);

FILL FILL_1__18778_ (
);

FILL FILL325280x247000 (
);

FILL FILL_1__18358_ (
);

AND2X2 _17636_ (
    .A(_6282__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [4]),
    .Y(_6558_)
);

OR2X2 _17216_ (
    .A(_6141_),
    .B(_6142_),
    .Y(_6143_)
);

NAND2X1 _12771_ (
    .A(_2330_),
    .B(_2335_),
    .Y(_2336_)
);

FILL FILL_0__12486_ (
);

OR2X2 _12351_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_1999_)
);

FILL FILL334400x49400 (
);

DFFSR _9978_ (
    .CLK(clk_bF$buf49),
    .D(_729_[6]),
    .Q(\datapath_1.regfile_1.regOut[12] [6]),
    .R(rst_bF$buf106),
    .S(vdd)
);

OR2X2 _9558_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_577_)
);

OR2X2 _9138_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_357_)
);

FILL FILL296400x123500 (
);

FILL FILL19760x276640 (
);

FILL FILL64600x251940 (
);

FILL FILL_0_BUFX2_insert580 (
);

FILL FILL3800x261820 (
);

FILL FILL_0_BUFX2_insert582 (
);

FILL FILL_0_BUFX2_insert584 (
);

OR2X2 _13976_ (
    .A(_3397_),
    .B(_3398_),
    .Y(_3399_)
);

FILL FILL_0_BUFX2_insert585 (
);

OR2X2 _13556_ (
    .A(ALUOut[22]),
    .B(_3079__bF$buf1),
    .Y(_3059_)
);

NOR2X1 _13136_ (
    .A(_2376__bF$buf2),
    .B(_2687_),
    .Y(_2688_)
);

FILL FILL_0_BUFX2_insert586 (
);

FILL FILL_0_BUFX2_insert587 (
);

FILL FILL_0_BUFX2_insert588 (
);

FILL FILL104120x340860 (
);

FILL FILL_0__14632_ (
);

FILL FILL_0__14212_ (
);

FILL FILL231040x64220 (
);

FILL FILL102600x187720 (
);

FILL FILL376960x276640 (
);

FILL FILL_0__15837_ (
);

OR2X2 _15702_ (
    .A(_4652_),
    .B(_4651_),
    .Y(_4653_)
);

FILL FILL_0__10972_ (
);

OR2X2 _18594_ (
    .A(_7500_),
    .B(_7497_),
    .Y(_7501_)
);

AND2X2 _18174_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_7088_)
);

FILL FILL_0__19250_ (
);

FILL FILL_1__12764_ (
);

AND2X2 _16907_ (
    .A(_4225__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_5839_)
);

FILL FILL13680x217360 (
);

FILL FILL_0__9771_ (
);

FILL FILL_0__11757_ (
);

OR2X2 _11622_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_1633_)
);

FILL FILL_0__11337_ (
);

OR2X2 _11202_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_1413_)
);

NOR2X1 _19379_ (
    .A(_6310__bF$buf1),
    .B(_8273_),
    .Y(_8274_)
);

AND2X2 _14094_ (
    .A(_3347__bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3500_)
);

DFFSR _8829_ (
    .CLK(clk_bF$buf52),
    .D(_135_[18]),
    .Q(\datapath_1.regfile_1.regOut[3] [18]),
    .R(rst_bF$buf55),
    .S(vdd)
);

BUFX2 _8409_ (
    .A(_1_[17]),
    .Y(memoryAddress[17])
);

FILL FILL_0__15590_ (
);

FILL FILL256120x256880 (
);

FILL FILL_0__15170_ (
);

FILL FILL343520x261820 (
);

FILL FILL_1__13969_ (
);

XNOR2X1 _12827_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2392_)
);

AND2X2 _12407_ (
    .A(_2036_),
    .B(_2035_),
    .Y(_1983_[26])
);

FILL FILL_1__14910_ (
);

FILL FILL273600x266760 (
);

AND2X2 _15299_ (
    .A(_4177__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_4256_)
);

FILL FILL_0__13903_ (
);

FILL FILL252320x88920 (
);

FILL FILL_1__17382_ (
);

AND2X2 _16660_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_5596_)
);

AND2X2 _16240_ (
    .A(_4167__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_5183_)
);

FILL FILL464360x74100 (
);

FILL FILL497800x103740 (
);

DFFSR _8582_ (
    .CLK(clk_bF$buf64),
    .D(_3_[29]),
    .Q(\datapath_1.regfile_1.regOut[1] [29]),
    .R(rst_bF$buf73),
    .S(vdd)
);

AND2X2 _17865_ (
    .A(_6783_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd1 [7])
);

FILL FILL491720x256880 (
);

AND2X2 _17445_ (
    .A(_6229__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_6370_)
);

OR2X2 _17025_ (
    .A(_5954_),
    .B(_5951_),
    .Y(_5955_)
);

AND2X2 _12580_ (
    .A(_2150_),
    .B(_2149_),
    .Y(_2143_[2])
);

OR2X2 _12160_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .B(_1916__bF$buf1),
    .Y(_1912_)
);

FILL FILL_0__18941_ (
);

FILL FILL_0__18521_ (
);

FILL FILL432440x242060 (
);

FILL FILL_0__18101_ (
);

OR2X2 _9787_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .B(_728__bF$buf3),
    .Y(_690_)
);

OR2X2 _9367_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_530__bF$buf2),
    .Y(_470_)
);

FILL FILL_0__8622_ (
);

FILL FILL_0__10608_ (
);

FILL FILL_1__14087_ (
);

FILL FILL238640x59280 (
);

OR2X2 _13785_ (
    .A(_3252_),
    .B(_3251_),
    .Y(_3253_)
);

AND2X2 _13365_ (
    .A(_2903_),
    .B(_2898_),
    .Y(_2904_)
);

FILL FILL468160x74100 (
);

FILL FILL_0__14021_ (
);

CLKBUF1 CLKBUF1_insert130 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf93)
);

CLKBUF1 CLKBUF1_insert131 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf92)
);

CLKBUF1 CLKBUF1_insert132 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf91)
);

CLKBUF1 CLKBUF1_insert133 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf90)
);

FILL FILL_0__9827_ (
);

CLKBUF1 CLKBUF1_insert134 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf89)
);

CLKBUF1 CLKBUF1_insert135 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf88)
);

CLKBUF1 CLKBUF1_insert136 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf87)
);

CLKBUF1 CLKBUF1_insert137 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf86)
);

CLKBUF1 CLKBUF1_insert138 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf85)
);

CLKBUF1 CLKBUF1_insert139 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf84)
);

FILL FILL408120x296400 (
);

AND2X2 _15931_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_4878_)
);

FILL FILL_0__15646_ (
);

OR2X2 _15511_ (
    .A(_4464_),
    .B(_4461_),
    .Y(_4465_)
);

FILL FILL_0__15226_ (
);

FILL FILL129960x187720 (
);

FILL FILL206720x133380 (
);

FILL FILL85120x207480 (
);

FILL FILL402800x29640 (
);

FILL FILL_1__17858_ (
);

FILL FILL266760x247000 (
);

OR2X2 _16716_ (
    .A(_5650_),
    .B(_5649_),
    .Y(_5651_)
);

FILL FILL_0__9580_ (
);

FILL FILL_0__11566_ (
);

OR2X2 _11851_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .B(_1784__bF$buf0),
    .Y(_1746_)
);

FILL FILL_0__9160_ (
);

OR2X2 _11431_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .B(_1586__bF$buf2),
    .Y(_1526_)
);

DFFSR _11011_ (
    .CLK(clk_bF$buf48),
    .D(_1257_[7]),
    .Q(\datapath_1.regfile_1.regOut[20] [7]),
    .R(rst_bF$buf21),
    .S(vdd)
);

OR2X2 _19188_ (
    .A(_8085_),
    .B(_8084_),
    .Y(_8086_)
);

FILL FILL487920x192660 (
);

OR2X2 _8638_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .B(_134__bF$buf3),
    .Y(_104_)
);

FILL FILL129200x311220 (
);

FILL FILL387600x286520 (
);

OR2X2 _12636_ (
    .A(_2200_),
    .B(_2188_),
    .Y(_2201_)
);

OR2X2 _12216_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_1929_)
);

FILL FILL310080x281580 (
);

FILL FILL301720x350740 (
);

FILL FILL47880x187720 (
);

FILL FILL_0__16184_ (
);

FILL FILL132240x251940 (
);

FILL FILL_1__15924_ (
);

FILL FILL502360x330980 (
);

FILL FILL_1__15504_ (
);

BUFX2 _8391_ (
    .A(_0_),
    .Y(MemWrite)
);

FILL FILL_0__14917_ (
);

FILL FILL47120x311220 (
);

FILL FILL326800x44460 (
);

AND2X2 _17674_ (
    .A(_6271__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_6595_)
);

OR2X2 _17254_ (
    .A(_6179_),
    .B(_6180_),
    .Y(_6181_)
);

FILL FILL_0__18750_ (
);

FILL FILL_0__18330_ (
);

DFFSR _9596_ (
    .CLK(clk_bF$buf83),
    .D(_531_[11]),
    .Q(\datapath_1.regfile_1.regOut[9] [11]),
    .R(rst_bF$buf17),
    .S(vdd)
);

AND2X2 _9176_ (
    .A(_382_),
    .B(_381_),
    .Y(_333_[24])
);

FILL FILL102600x4940 (
);

FILL FILL_0__8851_ (
);

FILL FILL_0__10417_ (
);

OR2X2 _10702_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .B(_1190__bF$buf1),
    .Y(_1160_)
);

AND2X2 _18879_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_7782_)
);

FILL FILL_0_BUFX2_insert960 (
);

AND2X2 _18459_ (
    .A(_6312__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_7368_)
);

FILL FILL230280x29640 (
);

FILL FILL_0_BUFX2_insert962 (
);

OR2X2 _18039_ (
    .A(_6951_),
    .B(_6954_),
    .Y(_6955_)
);

FILL FILL428640x39520 (
);

FILL FILL_0_BUFX2_insert964 (
);

FILL FILL_0_BUFX2_insert965 (
);

AND2X2 _13594_ (
    .A(ALUOp[0]),
    .B(PCSource[1]),
    .Y(_3089_)
);

XOR2X1 _13174_ (
    .A(_2718_),
    .B(_2449_),
    .Y(_2724_)
);

FILL FILL_0_BUFX2_insert966 (
);

FILL FILL_0_BUFX2_insert967 (
);

FILL FILL_0_BUFX2_insert968 (
);

AND2X2 _19400_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_8295_)
);

FILL FILL_0__19115_ (
);

FILL FILL_0__14670_ (
);

FILL FILL_0__14250_ (
);

FILL FILL293360x192660 (
);

FILL FILL_1__12629_ (
);

FILL FILL_0__9636_ (
);

DFFSR _11907_ (
    .CLK(clk_bF$buf105),
    .D(_1719_[0]),
    .Q(\datapath_1.regfile_1.regOut[27] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

OR2X2 _14799_ (
    .A(\datapath_1.rd2 [14]),
    .B(_3935__bF$buf1),
    .Y(_3899_)
);

OR2X2 _14379_ (
    .A(memoryOutData[3]),
    .B(_3737__bF$buf4),
    .Y(_3679_)
);

FILL FILL34200x44460 (
);

FILL FILL_0__15875_ (
);

AND2X2 _15740_ (
    .A(_4142__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_4690_)
);

FILL FILL_0__15455_ (
);

FILL FILL_0__15035_ (
);

OR2X2 _15320_ (
    .A(_4269_),
    .B(_4276_),
    .Y(_4277_)
);

FILL FILL98800x340860 (
);

FILL FILL_0__10590_ (
);

FILL FILL_0__10170_ (
);

FILL FILL_1__17247_ (
);

OR2X2 _10299_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_951_)
);

AND2X2 _16945_ (
    .A(_4183__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_5877_)
);

AND2X2 _16525_ (
    .A(_4160__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_5463_)
);

FILL FILL177840x44460 (
);

AND2X2 _16105_ (
    .A(_4228__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_5050_)
);

FILL FILL85120x345800 (
);

DFFSR _11660_ (
    .CLK(clk_bF$buf83),
    .D(_1587_[11]),
    .Q(\datapath_1.regfile_1.regOut[25] [11]),
    .R(rst_bF$buf17),
    .S(vdd)
);

AND2X2 _11240_ (
    .A(_1438_),
    .B(_1437_),
    .Y(_1389_[24])
);

FILL FILL373920x242060 (
);

AND2X2 _8867_ (
    .A(_216_),
    .B(_215_),
    .Y(_201_[7])
);

BUFX2 _8447_ (
    .A(_2_[23]),
    .Y(memoryWriteData[23])
);

FILL FILL381520x59280 (
);

FILL FILL411160x355680 (
);

FILL FILL_1__13587_ (
);

OR2X2 _12865_ (
    .A(_2429_),
    .B(_2415_),
    .Y(_2430_)
);

DFFSR _12445_ (
    .CLK(clk_bF$buf87),
    .D(_1983_[22]),
    .Q(\datapath_1.regfile_1.regOut[31] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

OR2X2 _12025_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .B(_1850__bF$buf4),
    .Y(_1842_)
);

FILL FILL_0__18806_ (
);

FILL FILL_0__13521_ (
);

FILL FILL110200x79040 (
);

FILL FILL_0__13101_ (
);

FILL FILL_1__9550_ (
);

FILL FILL_0__14306_ (
);

AND2X2 _17483_ (
    .A(_6229__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_6407_)
);

FILL FILL_0__17198_ (
);

OR2X2 _17063_ (
    .A(_5992_),
    .B(_5989_),
    .Y(_5993_)
);

FILL FILL495520x247000 (
);

FILL FILL_0_CLKBUF1_insert190 (
);

FILL FILL_0_CLKBUF1_insert192 (
);

FILL FILL_0_CLKBUF1_insert193 (
);

FILL FILL_0_CLKBUF1_insert194 (
);

FILL FILL_0_CLKBUF1_insert195 (
);

FILL FILL_0_CLKBUF1_insert196 (
);

FILL FILL_0__8660_ (
);

AND2X2 _10931_ (
    .A(_1272_),
    .B(_1271_),
    .Y(_1257_[7])
);

DFFSR _10511_ (
    .CLK(clk_bF$buf82),
    .D(_993_[23]),
    .Q(\datapath_1.regfile_1.regOut[16] [23]),
    .R(rst_bF$buf94),
    .S(vdd)
);

FILL FILL_0_CLKBUF1_insert198 (
);

FILL FILL_0__10226_ (
);

FILL FILL322240x306280 (
);

AND2X2 _18688_ (
    .A(_6317__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_7594_)
);

OR2X2 _18268_ (
    .A(_7178_),
    .B(_7179_),
    .Y(_7180_)
);

FILL FILL239400x316160 (
);

FILL FILL326800x321100 (
);

FILL FILL_0__19344_ (
);

FILL FILL_0_BUFX2_insert0 (
);

FILL FILL_0_BUFX2_insert1 (
);

FILL FILL_0_BUFX2_insert3 (
);

FILL FILL_0_BUFX2_insert5 (
);

OR2X2 _11716_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_1718__bF$buf3),
    .Y(_1676_)
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert9 (
);

OR2X2 _14188_ (
    .A(MemToReg_bF$buf0),
    .B(ALUOut[15]),
    .Y(_3570_)
);

FILL FILL_0__15684_ (
);

FILL FILL_1__17896_ (
);

FILL FILL_1__17476_ (
);

FILL FILL375440x212420 (
);

OR2X2 _16754_ (
    .A(_5688_),
    .B(_5687_),
    .Y(_5689_)
);

FILL FILL_0__16469_ (
);

FILL FILL_0__16049_ (
);

AND2X2 _16334_ (
    .A(_4208__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_5275_)
);

FILL FILL490960x83980 (
);

FILL FILL53200x14820 (
);

FILL FILL_0__17410_ (
);

OR2X2 _8676_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_129_)
);

FILL FILL430160x335920 (
);

FILL FILL304000x281580 (
);

OR2X2 _17959_ (
    .A(_6875_),
    .B(_6862_),
    .Y(_6876_)
);

OR2X2 _17539_ (
    .A(_6429_),
    .B(_6462_),
    .Y(_6463_)
);

OR2X2 _17119_ (
    .A(_6047_),
    .B(_6046_),
    .Y(_6048_)
);

FILL FILL_0__12389_ (
);

INVX1 _12674_ (
    .A(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2239_)
);

AND2X2 _12254_ (
    .A(_1954_),
    .B(_1953_),
    .Y(_1917_[18])
);

OR2X2 _18900_ (
    .A(_7799_),
    .B(_7802_),
    .Y(_7803_)
);

FILL FILL_0__18615_ (
);

FILL FILL_0__13750_ (
);

FILL FILL373160x286520 (
);

FILL FILL_0__13330_ (
);

FILL FILL209760x34580 (
);

FILL FILL196840x14820 (
);

OR2X2 _13879_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.mux_iord.din0 [21]),
    .Y(_3319_)
);

AND2X2 _13459_ (
    .A(_2991_),
    .B(_2905_),
    .Y(_2992_)
);

OR2X2 _13039_ (
    .A(_2387__bF$buf1),
    .B(_2596_),
    .Y(_2597_)
);

FILL FILL27360x143260 (
);

FILL FILL318440x108680 (
);

FILL FILL_0__14955_ (
);

OR2X2 _14820_ (
    .A(\datapath_1.rd2 [21]),
    .B(_3935__bF$buf3),
    .Y(_3913_)
);

FILL FILL_0__14535_ (
);

FILL FILL405840x113620 (
);

OR2X2 _14400_ (
    .A(memoryOutData[10]),
    .B(_3737__bF$buf1),
    .Y(_3693_)
);

FILL FILL459040x64220 (
);

INVX1 _17292_ (
    .A(\datapath_1.PCJump [26]),
    .Y(_6218_)
);

FILL FILL44840x153140 (
);

FILL FILL12920x365560 (
);

FILL FILL_1__16327_ (
);

FILL FILL_1__11882_ (
);

OR2X2 _15605_ (
    .A(_4556_),
    .B(_4557_),
    .Y(_4558_)
);

FILL FILL_0__10455_ (
);

OR2X2 _10740_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_1185_)
);

FILL FILL280440x316160 (
);

OR2X2 _10320_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_965_)
);

FILL FILL_0__10035_ (
);

FILL FILL422560x350740 (
);

AND2X2 _18497_ (
    .A(_6259__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_7406_)
);

AND2X2 _18077_ (
    .A(_6293__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_6992_)
);

FILL FILL16720x286520 (
);

FILL FILL288040x54340 (
);

FILL FILL_1__12247_ (
);

FILL FILL_0__9674_ (
);

AND2X2 _11945_ (
    .A(_1788_),
    .B(_1787_),
    .Y(_1785_[1])
);

DFFSR _11525_ (
    .CLK(clk_bF$buf29),
    .D(_1521_[5]),
    .Q(\datapath_1.regfile_1.regOut[24] [5]),
    .R(rst_bF$buf40),
    .S(vdd)
);

AND2X2 _11105_ (
    .A(_1368_),
    .B(_1367_),
    .Y(_1323_[22])
);

FILL FILL494000x113620 (
);

FILL FILL_0__12601_ (
);

FILL FILL_1__16080_ (
);

FILL FILL_0__15073_ (
);

FILL FILL452960x172900 (
);

FILL FILL388360x251940 (
);

FILL FILL_0__16698_ (
);

OR2X2 _16983_ (
    .A(_5910_),
    .B(_5913_),
    .Y(_5914_)
);

AND2X2 _16563_ (
    .A(_4230__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_5501_)
);

FILL FILL_0__16278_ (
);

OR2X2 _16143_ (
    .A(_5085_),
    .B(_5086_),
    .Y(_5087_)
);

OR2X2 _8485_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .B(_68__bF$buf2),
    .Y(_22_)
);

AND2X2 _17768_ (
    .A(_6297__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_6688_)
);

NOR3X1 _17348_ (
    .A(_6273_),
    .B(_6271__bF$buf0),
    .C(_6272__bF$buf1),
    .Y(_6274_)
);

FILL FILL_0__12198_ (
);

OR2X2 _12483_ (
    .A(_2074_),
    .B(_2065_),
    .Y(_2075_)
);

FILL FILL_1__19011_ (
);

DFFSR _12063_ (
    .CLK(clk_bF$buf14),
    .D(_1785_[27]),
    .Q(\datapath_1.regfile_1.regOut[28] [27]),
    .R(rst_bF$buf78),
    .S(vdd)
);

FILL FILL_0__18844_ (
);

FILL FILL435480x4940 (
);

FILL FILL145160x360620 (
);

FILL FILL411920x69160 (
);

FILL FILL259160x108680 (
);

FILL FILL_0__8525_ (
);

OR2X2 _13688_ (
    .A(_3169_),
    .B(_3166_),
    .Y(\datapath_1.mux_pcsrc.dout [13])
);

AOI21X1 _13268_ (
    .A(_2810_),
    .B(_2548_),
    .C(_2811_),
    .Y(_2812_)
);

FILL FILL_0__19209_ (
);

FILL FILL_0__14764_ (
);

FILL FILL46360x123500 (
);

FILL FILL_1__16976_ (
);

FILL FILL_0__15969_ (
);

AND2X2 _15834_ (
    .A(_4181__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [9]),
    .Y(_4783_)
);

FILL FILL_0__15549_ (
);

OR2X2 _15414_ (
    .A(_4366_),
    .B(_4369_),
    .Y(_4370_)
);

FILL FILL_0__10264_ (
);

FILL FILL498560x163020 (
);

FILL FILL248520x19760 (
);

FILL FILL_0__16910_ (
);

FILL FILL297920x370500 (
);

FILL FILL59280x4940 (
);

FILL FILL_0__19382_ (
);

FILL FILL206720x247000 (
);

OR2X2 _16619_ (
    .A(_5554_),
    .B(_5555_),
    .Y(_5556_)
);

FILL FILL_0__11469_ (
);

OR2X2 _11754_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_1701_)
);

FILL FILL_0__9063_ (
);

OR2X2 _11334_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_1481_)
);

FILL FILL_0__11049_ (
);

FILL FILL_0__12410_ (
);

FILL FILL145160x34580 (
);

AND2X2 _9902_ (
    .A(_746_),
    .B(_745_),
    .Y(_729_[8])
);

AOI21X1 _12959_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(_2364_),
    .C(_2365_),
    .Y(_2522_)
);

NOR3X1 _12539_ (
    .A(_2111_),
    .B(\control_1.op [0]),
    .C(\control_1.op [1]),
    .Y(_2128_)
);

AND2X2 _12119_ (
    .A(_1884_),
    .B(_1883_),
    .Y(_1851_[16])
);

FILL FILL_1_BUFX2_insert897 (
);

FILL FILL_1_BUFX2_insert899 (
);

OR2X2 _13900_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.PCJump [28]),
    .Y(_3333_)
);

FILL FILL_0__13615_ (
);

FILL FILL443080x306280 (
);

OR2X2 _16792_ (
    .A(_5725_),
    .B(_5718_),
    .Y(_5726_)
);

FILL FILL_0__16087_ (
);

AND2X2 _16372_ (
    .A(_4197__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_5313_)
);

FILL FILL_1__18299_ (
);

BUFX2 BUFX2_insert560 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf79)
);

BUFX2 BUFX2_insert561 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf78)
);

BUFX2 BUFX2_insert562 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf77)
);

BUFX2 BUFX2_insert563 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf76)
);

BUFX2 BUFX2_insert564 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf75)
);

AND2X2 _17997_ (
    .A(_6211__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_6913_)
);

BUFX2 BUFX2_insert565 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf74)
);

OR2X2 _17577_ (
    .A(_6496_),
    .B(_6499_),
    .Y(_6500_)
);

FILL FILL291080x217360 (
);

BUFX2 BUFX2_insert566 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf73)
);

AND2X2 _17157_ (
    .A(_4195__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_6085_)
);

BUFX2 BUFX2_insert567 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf72)
);

BUFX2 BUFX2_insert568 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf71)
);

BUFX2 BUFX2_insert569 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf70)
);

OR2X2 _12292_ (
    .A(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .B(_1982__bF$buf4),
    .Y(_1980_)
);

FILL FILL_1__19240_ (
);

FILL FILL22800x83980 (
);

FILL FILL_0__18233_ (
);

FILL FILL304000x217360 (
);

FILL FILL421800x133380 (
);

OR2X2 _9499_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .B(_596__bF$buf1),
    .Y(_538_)
);

DFFSR _9079_ (
    .CLK(clk_bF$buf108),
    .D(_267_[10]),
    .Q(\datapath_1.regfile_1.regOut[5] [10]),
    .R(rst_bF$buf56),
    .S(vdd)
);

FILL FILL_0__8754_ (
);

OR2X2 _10605_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_1115_)
);

FILL FILL_0_BUFX2_insert80 (
);

FILL FILL_0_BUFX2_insert82 (
);

FILL FILL_0_BUFX2_insert83 (
);

FILL FILL_0_BUFX2_insert84 (
);

FILL FILL_0_BUFX2_insert85 (
);

FILL FILL_0_BUFX2_insert86 (
);

AND2X2 _13497_ (
    .A(_3019_),
    .B(_3018_),
    .Y(_1_[2])
);

AND2X2 _13077_ (
    .A(_2632_),
    .B(_2630_),
    .Y(_2633_)
);

FILL FILL_0_BUFX2_insert88 (
);

FILL FILL_0__19438_ (
);

OR2X2 _19303_ (
    .A(_8198_),
    .B(_8194_),
    .Y(_8199_)
);

FILL FILL_0__14573_ (
);

FILL FILL456760x9880 (
);

FILL FILL_0__9119_ (
);

FILL FILL503880x163020 (
);

FILL FILL247760x153140 (
);

FILL FILL_1__16365_ (
);

FILL FILL430920x39520 (
);

FILL FILL287280x19760 (
);

AND2X2 _15643_ (
    .A(_4183__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_4595_)
);

NOR3X1 _15223_ (
    .A(_4140_),
    .B(\datapath_1.PCJump_22_bF$buf0 ),
    .C(_4153_),
    .Y(_4181_)
);

FILL FILL147440x247000 (
);

FILL FILL283480x232180 (
);

FILL FILL_0__19191_ (
);

OR2X2 _16848_ (
    .A(_5777_),
    .B(_5780_),
    .Y(_5781_)
);

AND2X2 _16428_ (
    .A(_4195__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_5368_)
);

OR2X2 _16008_ (
    .A(_4950_),
    .B(_4953_),
    .Y(_4954_)
);

OR2X2 _11983_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .B(_1850__bF$buf4),
    .Y(_1814_)
);

FILL FILL_0__9292_ (
);

OR2X2 _11563_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .B(_1652__bF$buf3),
    .Y(_1594_)
);

DFFSR _11143_ (
    .CLK(clk_bF$buf30),
    .D(_1323_[10]),
    .Q(\datapath_1.regfile_1.regOut[21] [10]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL439280x108680 (
);

FILL FILL494760x9880 (
);

FILL FILL_0__17924_ (
);

FILL FILL_0__17504_ (
);

FILL FILL163400x69160 (
);

FILL FILL438520x4940 (
);

FILL FILL318440x64220 (
);

FILL FILL335160x14820 (
);

OR2X2 _9711_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_659_)
);

INVX1 _12768_ (
    .A(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2333_)
);

OR2X2 _12348_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_1997_)
);

FILL FILL437760x276640 (
);

FILL FILL_0__18709_ (
);

FILL FILL109440x306280 (
);

FILL FILL_0__13844_ (
);

FILL FILL_0__13424_ (
);

FILL FILL_0__13004_ (
);

FILL FILL300200x247000 (
);

FILL FILL51680x271700 (
);

OR2X2 _16181_ (
    .A(_5123_),
    .B(_5124_),
    .Y(_5125_)
);

FILL FILL_1__9453_ (
);

FILL FILL366320x0 (
);

AND2X2 _14914_ (
    .A(_3955_),
    .B(_3954_),
    .Y(_3936_[9])
);

FILL FILL423320x103740 (
);

AND2X2 _17386_ (
    .A(_6249_),
    .B(\datapath_1.PCJump_27_bF$buf1 ),
    .Y(_6312_)
);

FILL FILL167200x69160 (
);

FILL FILL_0__18882_ (
);

FILL FILL_0__18462_ (
);

FILL FILL353400x108680 (
);

FILL FILL_1__11556_ (
);

FILL FILL27360x306280 (
);

FILL FILL_0__8983_ (
);

OR2X2 _10834_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .B(_1256__bF$buf1),
    .Y(_1228_)
);

FILL FILL_0__10549_ (
);

OR2X2 _10414_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .B(_1058__bF$buf4),
    .Y(_1008_)
);

FILL FILL418760x222300 (
);

DFFSR _19532_ (
    .CLK(clk_bF$buf55),
    .D(_8320_[9]),
    .Q(\datapath_1.regfile_1.regOut[0] [9]),
    .R(rst_bF$buf75),
    .S(vdd)
);

FILL FILL_0__19247_ (
);

AND2X2 _19112_ (
    .A(_6293__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_8011_)
);

FILL FILL_0__14382_ (
);

FILL FILL357200x350740 (
);

OR2X2 _11619_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_1631_)
);

FILL FILL_1__16594_ (
);

FILL FILL179360x128440 (
);

OR2X2 _15872_ (
    .A(_4818_),
    .B(_4819_),
    .Y(_4820_)
);

FILL FILL_0__15587_ (
);

OR2X2 _15452_ (
    .A(_4406_),
    .B(_4405_),
    .Y(_4407_)
);

FILL FILL_0__15167_ (
);

MUX2X1 _15032_ (
    .A(_4013_),
    .B(_4020_),
    .S(_4018_),
    .Y(_4021_)
);

FILL FILL11400x301340 (
);

FILL FILL228000x207480 (
);

AND2X2 _16657_ (
    .A(_4187__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_5593_)
);

AND2X2 _16237_ (
    .A(_4228__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_5180_)
);

DFFSR _11792_ (
    .CLK(clk_bF$buf98),
    .D(_1653_[14]),
    .Q(\datapath_1.regfile_1.regOut[26] [14]),
    .R(rst_bF$buf87),
    .S(vdd)
);

AND2X2 _11372_ (
    .A(_1506_),
    .B(_1505_),
    .Y(_1455_[25])
);

FILL FILL_0__11087_ (
);

FILL FILL_1__9509_ (
);

FILL FILL_0__17733_ (
);

FILL FILL_0__17313_ (
);

FILL FILL326800x281580 (
);

AND2X2 _8999_ (
    .A(_284_),
    .B(_283_),
    .Y(_267_[8])
);

DFFSR _8579_ (
    .CLK(clk_bF$buf54),
    .D(_3_[26]),
    .Q(\datapath_1.regfile_1.regOut[1] [26]),
    .R(rst_bF$buf14),
    .S(vdd)
);

FILL FILL_1__10827_ (
);

FILL FILL258400x163020 (
);

OR2X2 _9940_ (
    .A(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .B(_794__bF$buf2),
    .Y(_772_)
);

OR2X2 _9520_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .B(_596__bF$buf4),
    .Y(_552_)
);

DFFSR _9100_ (
    .CLK(clk_bF$buf9),
    .D(_267_[31]),
    .Q(\datapath_1.regfile_1.regOut[5] [31]),
    .R(rst_bF$buf23),
    .S(vdd)
);

AND2X2 _12997_ (
    .A(_2557_),
    .B(_2319_),
    .Y(_2558_)
);

AND2X2 _12577_ (
    .A(_2148_),
    .B(_2147_),
    .Y(_2143_[1])
);

FILL FILL_1__19105_ (
);

OR2X2 _12157_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .B(_1916__bF$buf1),
    .Y(_1910_)
);

FILL FILL163400x123500 (
);

FILL FILL78280x286520 (
);

OR2X2 _18803_ (
    .A(_7702_),
    .B(_7706_),
    .Y(_7707_)
);

FILL FILL_0__13653_ (
);

FILL FILL294120x242060 (
);

FILL FILL_0__8619_ (
);

FILL FILL459800x9880 (
);

BUFX2 BUFX2_insert1120 (
    .A(_1586_),
    .Y(_1586__bF$buf4)
);

BUFX2 BUFX2_insert1121 (
    .A(_1586_),
    .Y(_1586__bF$buf3)
);

BUFX2 BUFX2_insert1122 (
    .A(_1586_),
    .Y(_1586__bF$buf2)
);

BUFX2 BUFX2_insert1123 (
    .A(_1586_),
    .Y(_1586__bF$buf1)
);

BUFX2 BUFX2_insert1124 (
    .A(_1586_),
    .Y(_1586__bF$buf0)
);

BUFX2 BUFX2_insert1125 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf4 )
);

BUFX2 BUFX2_insert1126 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf3 )
);

BUFX2 BUFX2_insert1127 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf2 )
);

BUFX2 BUFX2_insert1128 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf1 )
);

FILL FILL_1__15445_ (
);

BUFX2 BUFX2_insert1129 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf0 )
);

FILL FILL_1__10580_ (
);

DFFSR _14723_ (
    .CLK(clk_bF$buf80),
    .D(_3804_[0]),
    .Q(\datapath_1.a [0]),
    .R(rst_bF$buf104),
    .S(vdd)
);

FILL FILL_0__14438_ (
);

FILL FILL_0__14018_ (
);

OR2X2 _14303_ (
    .A(vdd),
    .B(ALUOut[21]),
    .Y(_3648_)
);

FILL FILL313880x271700 (
);

BUFX2 BUFX2_insert940 (
    .A(_6287_),
    .Y(_6287__bF$buf2)
);

BUFX2 BUFX2_insert941 (
    .A(_6287_),
    .Y(_6287__bF$buf1)
);

BUFX2 BUFX2_insert942 (
    .A(_6287_),
    .Y(_6287__bF$buf0)
);

BUFX2 BUFX2_insert943 (
    .A(_1058_),
    .Y(_1058__bF$buf4)
);

BUFX2 BUFX2_insert944 (
    .A(_1058_),
    .Y(_1058__bF$buf3)
);

BUFX2 BUFX2_insert945 (
    .A(_1058_),
    .Y(_1058__bF$buf2)
);

BUFX2 BUFX2_insert946 (
    .A(_1058_),
    .Y(_1058__bF$buf1)
);

OR2X2 _17195_ (
    .A(_6121_),
    .B(_6122_),
    .Y(_6123_)
);

BUFX2 BUFX2_insert947 (
    .A(_1058_),
    .Y(_1058__bF$buf0)
);

BUFX2 BUFX2_insert948 (
    .A(_4065_),
    .Y(_4065__bF$buf7)
);

FILL FILL357200x49400 (
);

BUFX2 BUFX2_insert949 (
    .A(_4065_),
    .Y(_4065__bF$buf6)
);

FILL FILL_0__18691_ (
);

OR2X2 _15928_ (
    .A(_4875_),
    .B(_4860_),
    .Y(_4876_)
);

AND2X2 _15508_ (
    .A(_4236__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_4462_)
);

FILL FILL_0__8792_ (
);

FILL FILL_0__10778_ (
);

FILL FILL_0__10358_ (
);

DFFSR _10643_ (
    .CLK(clk_bF$buf55),
    .D(_1059_[26]),
    .Q(\datapath_1.regfile_1.regOut[17] [26]),
    .R(rst_bF$buf27),
    .S(vdd)
);

AND2X2 _10223_ (
    .A(_920_),
    .B(_919_),
    .Y(_861_[29])
);

FILL FILL406600x59280 (
);

FILL FILL_0__19476_ (
);

FILL FILL_0__19056_ (
);

OR2X2 _19341_ (
    .A(_8236_),
    .B(_8229_),
    .Y(_8237_)
);

FILL FILL_0__14191_ (
);

FILL FILL_0__9577_ (
);

OR2X2 _11848_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .B(_1784__bF$buf3),
    .Y(_1744_)
);

OR2X2 _11428_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .B(_1586__bF$buf0),
    .Y(_1524_)
);

DFFSR _11008_ (
    .CLK(clk_bF$buf73),
    .D(_1257_[4]),
    .Q(\datapath_1.regfile_1.regOut[20] [4]),
    .R(rst_bF$buf39),
    .S(vdd)
);

FILL FILL_1__13511_ (
);

FILL FILL123120x256880 (
);

FILL FILL279680x172900 (
);

FILL FILL484880x350740 (
);

FILL FILL_0__15396_ (
);

OR2X2 _15681_ (
    .A(_4628_),
    .B(_4631_),
    .Y(_4632_)
);

OR2X2 _15261_ (
    .A(_4215_),
    .B(_4218_),
    .Y(_4219_)
);

FILL FILL15960x217360 (
);

FILL FILL_0__13709_ (
);

FILL FILL118560x375440 (
);

OR2X2 _16886_ (
    .A(_5815_),
    .B(_5818_),
    .Y(_5819_)
);

AND2X2 _16466_ (
    .A(_4154__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_5405_)
);

OR2X2 _16046_ (
    .A(_4990_),
    .B(_4991_),
    .Y(_4992_)
);

OR2X2 _11181_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_1399_)
);

FILL FILL_0__17962_ (
);

FILL FILL258400x256880 (
);

FILL FILL41040x256880 (
);

FILL FILL_1__10216_ (
);

FILL FILL45600x271700 (
);

AND2X2 _12386_ (
    .A(_2022_),
    .B(_2021_),
    .Y(_1983_[19])
);

FILL FILL104120x202540 (
);

FILL FILL_0__18747_ (
);

AND2X2 _18612_ (
    .A(_6259__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_7519_)
);

FILL FILL_0__18327_ (
);

FILL FILL_0__13462_ (
);

FILL FILL_0__13042_ (
);

FILL FILL362520x177840 (
);

FILL FILL234080x59280 (
);

FILL FILL_0__8428_ (
);

FILL FILL158840x335920 (
);

FILL FILL216600x118560 (
);

FILL FILL_0__14667_ (
);

OR2X2 _14952_ (
    .A(\datapath_1.mux_pcsrc.dout [22]),
    .B(_4001__bF$buf2),
    .Y(_3981_)
);

OR2X2 _14532_ (
    .A(memoryOutData[11]),
    .B(_3803__bF$buf3),
    .Y(_3761_)
);

OR2X2 _14112_ (
    .A(_3515_),
    .B(_3514_),
    .Y(_3516_)
);

FILL FILL357960x296400 (
);

FILL FILL_0__18080_ (
);

FILL FILL61560x19760 (
);

FILL FILL_1__16459_ (
);

OR2X2 _15737_ (
    .A(_4687_),
    .B(_4656_),
    .Y(_4688_)
);

AND2X2 _15317_ (
    .A(_4208__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_4274_)
);

OR2X2 _10872_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_1253_)
);

FILL FILL_0__10587_ (
);

OR2X2 _10452_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_1033_)
);

FILL FILL_0__10167_ (
);

OR2X2 _10032_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_813_)
);

BUFX2 BUFX2_insert90 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf4 )
);

BUFX2 BUFX2_insert91 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf3 )
);

BUFX2 BUFX2_insert92 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf2 )
);

BUFX2 BUFX2_insert93 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf1 )
);

BUFX2 BUFX2_insert94 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf0 )
);

BUFX2 BUFX2_insert95 (
    .A(_4208_),
    .Y(_4208__bF$buf4)
);

BUFX2 BUFX2_insert96 (
    .A(_4208_),
    .Y(_4208__bF$buf3)
);

BUFX2 BUFX2_insert97 (
    .A(_4208_),
    .Y(_4208__bF$buf2)
);

BUFX2 BUFX2_insert98 (
    .A(_4208_),
    .Y(_4208__bF$buf1)
);

BUFX2 BUFX2_insert99 (
    .A(_4208_),
    .Y(_4208__bF$buf0)
);

FILL FILL_0__19285_ (
);

AND2X2 _19150_ (
    .A(_6289__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_8049_)
);

FILL FILL343520x123500 (
);

AND2X2 _8600_ (
    .A(_78_),
    .B(_77_),
    .Y(_69_[4])
);

FILL FILL17480x321100 (
);

FILL FILL_0__9386_ (
);

DFFSR _11657_ (
    .CLK(clk_bF$buf22),
    .D(_1587_[8]),
    .Q(\datapath_1.regfile_1.regOut[25] [8]),
    .R(rst_bF$buf7),
    .S(vdd)
);

FILL FILL_1__18605_ (
);

AND2X2 _11237_ (
    .A(_1436_),
    .B(_1435_),
    .Y(_1389_[23])
);

FILL FILL_0__12733_ (
);

FILL FILL250800x19760 (
);

AND2X2 _15490_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_4444_)
);

AND2X2 _15070_ (
    .A(_4057_),
    .B(_4041_),
    .Y(_4058_)
);

FILL FILL65360x19760 (
);

OR2X2 _9805_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .B(_728__bF$buf0),
    .Y(_702_)
);

FILL FILL87400x207480 (
);

FILL FILL_1__14945_ (
);

FILL FILL478800x123500 (
);

FILL FILL_0__13938_ (
);

FILL FILL_0__13518_ (
);

OR2X2 _13803_ (
    .A(_3266_),
    .B(_3267_),
    .Y(_3268_)
);

OR2X2 _16695_ (
    .A(_5630_),
    .B(_5623_),
    .Y(_5631_)
);

OR2X2 _16275_ (
    .A(_5216_),
    .B(_5215_),
    .Y(_5217_)
);

FILL FILL345800x44460 (
);

FILL FILL_0__17351_ (
);

FILL FILL_1__10025_ (
);

FILL FILL231040x217360 (
);

DFFSR _12195_ (
    .CLK(clk_bF$buf30),
    .D(_1851_[30]),
    .Q(\datapath_1.regfile_1.regOut[29] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL229520x291460 (
);

FILL FILL_0__18976_ (
);

FILL FILL_0__18556_ (
);

AND2X2 _18841_ (
    .A(_6244__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_7744_)
);

OR2X2 _18421_ (
    .A(_7329_),
    .B(_7330_),
    .Y(_7331_)
);

OR2X2 _18001_ (
    .A(_6915_),
    .B(_6916_),
    .Y(_6917_)
);

FILL FILL_0__13691_ (
);

FILL FILL_0__8657_ (
);

AND2X2 _10928_ (
    .A(_1270_),
    .B(_1269_),
    .Y(_1257_[6])
);

DFFSR _10508_ (
    .CLK(clk_bF$buf100),
    .D(_993_[20]),
    .Q(\datapath_1.regfile_1.regOut[16] [20]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL504640x330980 (
);

FILL FILL_1__15483_ (
);

FILL FILL_1__15063_ (
);

FILL FILL349600x44460 (
);

AND2X2 _19206_ (
    .A(_6238__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_8104_)
);

FILL FILL_0__14896_ (
);

AND2X2 _14761_ (
    .A(_3873_),
    .B(_3872_),
    .Y(_3870_[1])
);

FILL FILL_0__14056_ (
);

DFFSR _14341_ (
    .CLK(clk_bF$buf20),
    .D(_3606_[5]),
    .Q(ALUOut[5]),
    .R(rst_bF$buf29),
    .S(vdd)
);

FILL FILL453720x222300 (
);

FILL FILL276640x29640 (
);

FILL FILL460560x29640 (
);

FILL FILL142880x365560 (
);

FILL FILL330600x4940 (
);

FILL FILL392160x158080 (
);

FILL FILL389120x301340 (
);

AND2X2 _15966_ (
    .A(_4172__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_4913_)
);

AND2X2 _15546_ (
    .A(_4499_),
    .B(_4065__bF$buf0),
    .Y(\datapath_1.rd2 [4])
);

AND2X2 _15126_ (
    .A(_4100_),
    .B(_4102_),
    .Y(_4103_)
);

FILL FILL_0__10396_ (
);

OR2X2 _10681_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .B(_1190__bF$buf1),
    .Y(_1146_)
);

DFFSR _10261_ (
    .CLK(clk_bF$buf71),
    .D(_861_[31]),
    .Q(\datapath_1.regfile_1.regOut[14] [31]),
    .R(rst_bF$buf35),
    .S(vdd)
);

FILL FILL_0__16202_ (
);

FILL FILL470440x138320 (
);

FILL FILL240920x242060 (
);

OR2X2 _11886_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_1769_)
);

FILL FILL_0__9195_ (
);

OR2X2 _11466_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_1549_)
);

OR2X2 _11046_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_1329_)
);

FILL FILL_0__17827_ (
);

FILL FILL_0__12962_ (
);

FILL FILL_0__12542_ (
);

FILL FILL_0__12122_ (
);

FILL FILL310840x103740 (
);

DFFSR _9614_ (
    .CLK(clk_bF$buf5),
    .D(_531_[29]),
    .Q(\datapath_1.regfile_1.regOut[9] [29]),
    .R(rst_bF$buf37),
    .S(vdd)
);

FILL FILL_1__8991_ (
);

FILL FILL_1__14334_ (
);

AND2X2 _13612_ (
    .A(_3081__bF$buf3),
    .B(ALUOut[3]),
    .Y(_3104_)
);

FILL FILL384560x44460 (
);

FILL FILL87400x345800 (
);

FILL FILL218880x217360 (
);

AND2X2 _16084_ (
    .A(_4172__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_5029_)
);

FILL FILL177080x44460 (
);

FILL FILL413440x355680 (
);

FILL FILL_0__17580_ (
);

FILL FILL_1__15959_ (
);

OR2X2 _14817_ (
    .A(\datapath_1.rd2 [20]),
    .B(_3935__bF$buf3),
    .Y(_3911_)
);

FILL FILL430920x365560 (
);

FILL FILL_1__16900_ (
);

FILL FILL500080x266760 (
);

FILL FILL427880x316160 (
);

AND2X2 _17289_ (
    .A(_6204_),
    .B(_6214_),
    .Y(_6215_)
);

AND2X2 _18650_ (
    .A(_6289__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_7556_)
);

FILL FILL_0__18365_ (
);

OR2X2 _18230_ (
    .A(_7141_),
    .B(_7142_),
    .Y(_7143_)
);

FILL FILL_0__13080_ (
);

FILL FILL_0__8886_ (
);

FILL FILL_0__8466_ (
);

OR2X2 _10737_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_1183_)
);

OR2X2 _10317_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_963_)
);

FILL FILL_1__12400_ (
);

FILL FILL_0__11813_ (
);

AND2X2 _19435_ (
    .A(_8325_),
    .B(_8324_),
    .Y(_8320_[2])
);

OR2X2 _19015_ (
    .A(_7915_),
    .B(_7908_),
    .Y(_7916_)
);

DFFSR _14990_ (
    .CLK(clk_bF$buf50),
    .D(_3936_[9]),
    .Q(\datapath_1.mux_iord.din0 [9]),
    .R(rst_bF$buf86),
    .S(vdd)
);

FILL FILL_0__14285_ (
);

OR2X2 _14570_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump [26]),
    .Y(_3786_)
);

OR2X2 _14150_ (
    .A(\datapath_1.Data [2]),
    .B(_3605__bF$buf1),
    .Y(_3545_)
);

FILL FILL379240x256880 (
);

FILL FILL135280x74100 (
);

OR2X2 _15775_ (
    .A(_4723_),
    .B(_4724_),
    .Y(_4725_)
);

AND2X2 _15355_ (
    .A(_4187__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_4311_)
);

DFFSR _10490_ (
    .CLK(clk_bF$buf56),
    .D(_993_[2]),
    .Q(\datapath_1.regfile_1.regOut[16] [2]),
    .R(rst_bF$buf30),
    .S(vdd)
);

AND2X2 _10070_ (
    .A(_838_),
    .B(_837_),
    .Y(_795_[21])
);

FILL FILL310840x330980 (
);

FILL FILL_0__16851_ (
);

FILL FILL_0__16431_ (
);

OR2X2 _11695_ (
    .A(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .B(_1718__bF$buf0),
    .Y(_1662_)
);

FILL FILL_1__18223_ (
);

DFFSR _11275_ (
    .CLK(clk_bF$buf13),
    .D(_1389_[13]),
    .Q(\datapath_1.regfile_1.regOut[22] [13]),
    .R(rst_bF$buf90),
    .S(vdd)
);

OR2X2 _17921_ (
    .A(_6837_),
    .B(_6838_),
    .Y(_6839_)
);

FILL FILL_0__17216_ (
);

AND2X2 _17501_ (
    .A(_6264__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_6425_)
);

FILL FILL_0__12771_ (
);

FILL FILL_0__12351_ (
);

DFFSR _9843_ (
    .CLK(clk_bF$buf96),
    .D(_663_[0]),
    .Q(\datapath_1.regfile_1.regOut[11] [0]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9423_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_507_)
);

OR2X2 _9003_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_287_)
);

OR2X2 _18706_ (
    .A(_7604_),
    .B(_7611_),
    .Y(_7612_)
);

OR2X2 _13841_ (
    .A(\datapath_1.a [8]),
    .B(_3342__bF$buf4),
    .Y(_3294_)
);

FILL FILL_0__13556_ (
);

FILL FILL192280x14820 (
);

FILL FILL_0__13136_ (
);

AND2X2 _13421_ (
    .A(_2952_),
    .B(_2955_),
    .Y(_2956_)
);

INVX1 _13001_ (
    .A(_2561_),
    .Y(\datapath_1.ALUResult [27])
);

FILL FILL432440x335920 (
);

OR2X2 _14626_ (
    .A(\datapath_1.a [0]),
    .B(vdd),
    .Y(_3868_)
);

OR2X2 _14206_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[21]),
    .Y(_3582_)
);

AND2X2 _17098_ (
    .A(_4217__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_6027_)
);

FILL FILL_0__15702_ (
);

FILL FILL367840x98800 (
);

FILL FILL_0__18174_ (
);

FILL FILL_1__11688_ (
);

OR2X2 _10966_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .B(_1322__bF$buf3),
    .Y(_1296_)
);

OR2X2 _10546_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .B(_1124__bF$buf0),
    .Y(_1076_)
);

DFFSR _10126_ (
    .CLK(clk_bF$buf60),
    .D(_795_[25]),
    .Q(\datapath_1.regfile_1.regOut[13] [25]),
    .R(rst_bF$buf101),
    .S(vdd)
);

FILL FILL_0__16907_ (
);

FILL FILL29640x143260 (
);

FILL FILL243200x74100 (
);

FILL FILL_0__11622_ (
);

OR2X2 _19244_ (
    .A(_8137_),
    .B(_8140_),
    .Y(_8141_)
);

FILL FILL_0__14094_ (
);

FILL FILL145920x256880 (
);

FILL FILL_1__13834_ (
);

FILL FILL_0__12827_ (
);

FILL FILL_0__12407_ (
);

FILL FILL232560x167960 (
);

OR2X2 _15584_ (
    .A(_4533_),
    .B(_4536_),
    .Y(_4537_)
);

NOR3X1 _15164_ (
    .A(_4125_),
    .B(_4059_),
    .C(_4011_),
    .Y(\datapath_1.regfile_1.regEn [28])
);

FILL FILL_1__8436_ (
);

FILL FILL450680x291460 (
);

FILL FILL471200x24700 (
);

FILL FILL201400x59280 (
);

FILL FILL69920x103740 (
);

AND2X2 _16789_ (
    .A(_4208__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_5723_)
);

AND2X2 _16369_ (
    .A(_4200__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_5310_)
);

FILL FILL_1__18872_ (
);

AND2X2 _11084_ (
    .A(_1354_),
    .B(_1353_),
    .Y(_1323_[15])
);

FILL FILL_0__17865_ (
);

FILL FILL373160x148200 (
);

FILL FILL_0__17445_ (
);

OR2X2 _17730_ (
    .A(_6647_),
    .B(_6650_),
    .Y(_6651_)
);

FILL FILL_0__17025_ (
);

AND2X2 _17310_ (
    .A(_6235_),
    .B(\datapath_1.PCJump_27_bF$buf0 ),
    .Y(_6236_)
);

FILL FILL63840x256880 (
);

FILL FILL386840x330980 (
);

FILL FILL_0__12580_ (
);

FILL FILL_0__12160_ (
);

FILL FILL_1__10959_ (
);

OR2X2 _9652_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .B(_662__bF$buf2),
    .Y(_620_)
);

OR2X2 _9232_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(_464__bF$buf0),
    .Y(_400_)
);

FILL FILL203680x54340 (
);

OR2X2 _12289_ (
    .A(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .B(_1982__bF$buf1),
    .Y(_1978_)
);

AND2X2 _18935_ (
    .A(_6282__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_7837_)
);

AND2X2 _18515_ (
    .A(_7423_),
    .B(_4065__bF$buf3),
    .Y(\datapath_1.rd1 [17])
);

FILL FILL503120x291460 (
);

FILL FILL_0__13785_ (
);

AND2X2 _13650_ (
    .A(_3087__bF$buf1),
    .B(\datapath_1.ALUResult [8]),
    .Y(_3137_)
);

FILL FILL247000x281580 (
);

AND2X2 _13230_ (
    .A(_2776_),
    .B(_2772_),
    .Y(_2777_)
);

FILL FILL_1__15577_ (
);

DFFSR _14855_ (
    .CLK(clk_bF$buf38),
    .D(_3870_[3]),
    .Q(_2_[3]),
    .R(rst_bF$buf70),
    .S(vdd)
);

OR2X2 _14435_ (
    .A(vdd),
    .B(\datapath_1.Data [22]),
    .Y(_3716_)
);

OR2X2 _14015_ (
    .A(_3432_),
    .B(_3429_),
    .Y(\datapath_1.alu_1.ALUInB [13])
);

FILL FILL_0__15931_ (
);

FILL FILL_0__15511_ (
);

FILL FILL_1__11077_ (
);

FILL FILL_1__17723_ (
);

DFFSR _10775_ (
    .CLK(clk_bF$buf76),
    .D(_1125_[29]),
    .Q(\datapath_1.regfile_1.regOut[18] [29]),
    .R(rst_bF$buf110),
    .S(vdd)
);

AND2X2 _10355_ (
    .A(_988_),
    .B(_987_),
    .Y(_927_[30])
);

FILL FILL_0__16716_ (
);

FILL FILL48640x123500 (
);

FILL FILL_0__11851_ (
);

FILL FILL_0__19188_ (
);

OR2X2 _19473_ (
    .A(gnd),
    .B(_8385__bF$buf3),
    .Y(_8351_)
);

AND2X2 _19053_ (
    .A(_6211__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_7953_)
);

OR2X2 _8923_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .B(_266__bF$buf3),
    .Y(_254_)
);

OR2X2 _8503_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .B(_68__bF$buf2),
    .Y(_34_)
);

OR2X2 _12921_ (
    .A(_2485_),
    .B(_2484_),
    .Y(_2486_)
);

FILL FILL_0__12636_ (
);

FILL FILL_0__12216_ (
);

XOR2X1 _12501_ (
    .A(\control_1.reg_state.dout [2]),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2099_)
);

FILL FILL_1_BUFX2_insert517 (
);

FILL FILL_1_BUFX2_insert519 (
);

AND2X2 _15393_ (
    .A(_4135__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .Y(_4349_)
);

OR2X2 _9708_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_657_)
);

FILL FILL141360x301340 (
);

FILL FILL299440x276640 (
);

AND2X2 _13706_ (
    .A(_3087__bF$buf2),
    .B(\datapath_1.ALUResult [16]),
    .Y(_3185_)
);

FILL FILL375440x34580 (
);

OR2X2 _16598_ (
    .A(_5534_),
    .B(_5533_),
    .Y(_5535_)
);

OR2X2 _16178_ (
    .A(_5121_),
    .B(_5120_),
    .Y(_5122_)
);

FILL FILL_0__17674_ (
);

FILL FILL41800x83980 (
);

FILL FILL17480x281580 (
);

AND2X2 _9881_ (
    .A(_732_),
    .B(_731_),
    .Y(_729_[1])
);

DFFSR _9461_ (
    .CLK(clk_bF$buf104),
    .D(_465_[5]),
    .Q(\datapath_1.regfile_1.regOut[8] [5]),
    .R(rst_bF$buf80),
    .S(vdd)
);

AND2X2 _9041_ (
    .A(_312_),
    .B(_311_),
    .Y(_267_[22])
);

AND2X2 _12098_ (
    .A(_1870_),
    .B(_1869_),
    .Y(_1851_[9])
);

FILL FILL_1__19046_ (
);

FILL FILL_0__10702_ (
);

FILL FILL_0__18879_ (
);

OR2X2 _18744_ (
    .A(_7648_),
    .B(_7647_),
    .Y(_7649_)
);

AND2X2 _18324_ (
    .A(_6206__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_7235_)
);

FILL FILL_0__18039_ (
);

FILL FILL_0__13594_ (
);

FILL FILL_0__13174_ (
);

FILL FILL431680x330980 (
);

FILL FILL257640x138320 (
);

FILL FILL_0__9921_ (
);

FILL FILL_0__9501_ (
);

DFFSR _19529_ (
    .CLK(clk_bF$buf70),
    .D(_8320_[6]),
    .Q(\datapath_1.regfile_1.regOut[0] [6]),
    .R(rst_bF$buf66),
    .S(vdd)
);

AND2X2 _19109_ (
    .A(_6328__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_8008_)
);

FILL FILL293360x217360 (
);

FILL FILL_0__14799_ (
);

OR2X2 _14664_ (
    .A(\datapath_1.rd1 [12]),
    .B(_3869__bF$buf4),
    .Y(_3829_)
);

OR2X2 _14244_ (
    .A(\datapath_1.ALUResult [1]),
    .B(_3671__bF$buf4),
    .Y(_3609_)
);

FILL FILL_0__15320_ (
);

FILL FILL335160x345800 (
);

OR2X2 _15869_ (
    .A(_4816_),
    .B(_4815_),
    .Y(_4817_)
);

OR2X2 _15449_ (
    .A(_4403_),
    .B(_4388_),
    .Y(_4404_)
);

NOR2X1 _15029_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_4018_)
);

OR2X2 _10584_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_1101_)
);

FILL FILL_0__10299_ (
);

FILL FILL417240x49400 (
);

FILL FILL_1__17112_ (
);

OR2X2 _10164_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_881_)
);

FILL FILL_0__16945_ (
);

FILL FILL_0__16525_ (
);

AND2X2 _16810_ (
    .A(_4225__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_5744_)
);

FILL FILL_0__11240_ (
);

OR2X2 _19282_ (
    .A(_8178_),
    .B(_8177_),
    .Y(_8179_)
);

FILL FILL332880x143260 (
);

AND2X2 _8732_ (
    .A(_146_),
    .B(_145_),
    .Y(_135_[5])
);

FILL FILL_1__18737_ (
);

DFFSR _11789_ (
    .CLK(clk_bF$buf79),
    .D(_1653_[11]),
    .Q(\datapath_1.regfile_1.regOut[26] [11]),
    .R(rst_bF$buf57),
    .S(vdd)
);

AND2X2 _11369_ (
    .A(_1504_),
    .B(_1503_),
    .Y(_1455_[24])
);

FILL FILL_1__13452_ (
);

OR2X2 _12730_ (
    .A(_2289_),
    .B(_2294_),
    .Y(_2295_)
);

DFFSR _12310_ (
    .CLK(clk_bF$buf78),
    .D(_1917_[16]),
    .Q(\datapath_1.regfile_1.regOut[30] [16]),
    .R(rst_bF$buf110),
    .S(vdd)
);

FILL FILL131480x256880 (
);

OR2X2 _9937_ (
    .A(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .B(_794__bF$buf4),
    .Y(_770_)
);

OR2X2 _9517_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .B(_596__bF$buf0),
    .Y(_550_)
);

FILL FILL304760x276640 (
);

AND2X2 _13935_ (
    .A(_3350__bF$buf0),
    .B(_2_[2]),
    .Y(_3364_)
);

AND2X2 _13515_ (
    .A(_3031_),
    .B(_3030_),
    .Y(_1_[8])
);

FILL FILL129200x133380 (
);

BUFX2 BUFX2_insert1090 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf4 )
);

BUFX2 BUFX2_insert1091 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf3 )
);

BUFX2 BUFX2_insert1092 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf2 )
);

FILL FILL_0__17483_ (
);

FILL FILL55480x103740 (
);

FILL FILL186200x69160 (
);

FILL FILL_0__17063_ (
);

BUFX2 BUFX2_insert1093 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf1 )
);

BUFX2 BUFX2_insert1094 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf0 )
);

BUFX2 BUFX2_insert1095 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf4 )
);

BUFX2 BUFX2_insert1096 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf3 )
);

BUFX2 BUFX2_insert1097 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf2 )
);

BUFX2 BUFX2_insert1098 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf1 )
);

BUFX2 BUFX2_insert1099 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf0 )
);

FILL FILL36480x261820 (
);

OR2X2 _9690_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_645_)
);

OR2X2 _9270_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_425_)
);

FILL FILL_1_CLKBUF1_insert223 (
);

FILL FILL268280x49400 (
);

FILL FILL_0__10931_ (
);

OR2X2 _18973_ (
    .A(_7872_),
    .B(_7873_),
    .Y(_7874_)
);

OR2X2 _18553_ (
    .A(_7460_),
    .B(_7457_),
    .Y(_7461_)
);

FILL FILL_0__18268_ (
);

AND2X2 _18133_ (
    .A(_6300__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_7047_)
);

FILL FILL201400x266760 (
);

FILL FILL224200x350740 (
);

FILL FILL_0__9310_ (
);

FILL FILL364800x133380 (
);

AND2X2 _19338_ (
    .A(_6232__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_8234_)
);

FILL FILL70680x187720 (
);

AND2X2 _14893_ (
    .A(_3941_),
    .B(_3940_),
    .Y(_3936_[2])
);

DFFSR _14473_ (
    .CLK(clk_bF$buf23),
    .D(_3672_[8]),
    .Q(\datapath_1.Data [8]),
    .R(rst_bF$buf33),
    .S(vdd)
);

OR2X2 _14053_ (
    .A(_3463_),
    .B(_3464_),
    .Y(_3465_)
);

FILL FILL_1__13928_ (
);

FILL FILL3800x153140 (
);

FILL FILL416480x207480 (
);

FILL FILL503880x212420 (
);

AND2X2 _15678_ (
    .A(_4230__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_4629_)
);

NOR3X1 _15258_ (
    .A(_4126_),
    .B(\datapath_1.PCJump [18]),
    .C(_4153_),
    .Y(_4216_)
);

OR2X2 _10393_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(_1058__bF$buf3),
    .Y(_994_)
);

FILL FILL_1__17341_ (
);

FILL FILL_0__16334_ (
);

FILL FILL423320x177840 (
);

OR2X2 _19091_ (
    .A(_7989_),
    .B(_7990_),
    .Y(_7991_)
);

DFFSR _8961_ (
    .CLK(clk_bF$buf34),
    .D(_201_[21]),
    .Q(\datapath_1.regfile_1.regOut[4] [21]),
    .R(rst_bF$buf71),
    .S(vdd)
);

OR2X2 _8541_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_59_)
);

FILL FILL437760x138320 (
);

FILL FILL_1__18546_ (
);

OR2X2 _11598_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_1617_)
);

OR2X2 _11178_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_1397_)
);

FILL FILL_0__17539_ (
);

OR2X2 _17824_ (
    .A(_6741_),
    .B(_6742_),
    .Y(_6743_)
);

OR2X2 _17404_ (
    .A(_6327_),
    .B(_6329_),
    .Y(_6330_)
);

FILL FILL_0__17119_ (
);

FILL FILL_0__12674_ (
);

OR2X2 _9746_ (
    .A(\datapath_1.regfile_1.regOut[11] [0]),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .Y(_727_)
);

AND2X2 _9326_ (
    .A(_462_),
    .B(_461_),
    .Y(_399_[31])
);

FILL FILL268280x360620 (
);

FILL FILL161120x242060 (
);

FILL FILL_1__14886_ (
);

OR2X2 _18609_ (
    .A(_7508_),
    .B(_7515_),
    .Y(_7516_)
);

FILL FILL_0__13879_ (
);

FILL FILL_0__13459_ (
);

OR2X2 _13744_ (
    .A(_3217_),
    .B(_3214_),
    .Y(\datapath_1.mux_pcsrc.dout [21])
);

OR2X2 _13324_ (
    .A(_2157__bF$buf1),
    .B(_2864_),
    .Y(_2865_)
);

FILL FILL_0__17292_ (
);

OR2X2 _14949_ (
    .A(\datapath_1.mux_pcsrc.dout [21]),
    .B(_4001__bF$buf1),
    .Y(_3979_)
);

OR2X2 _14529_ (
    .A(memoryOutData[10]),
    .B(_3803__bF$buf0),
    .Y(_3759_)
);

OR2X2 _14109_ (
    .A(_3511_),
    .B(_3512_),
    .Y(_3513_)
);

FILL FILL440040x202540 (
);

FILL FILL405840x44460 (
);

FILL FILL_1__19084_ (
);

FILL FILL_0__10740_ (
);

FILL FILL296400x242060 (
);

FILL FILL_0__10320_ (
);

OR2X2 _18782_ (
    .A(_7682_),
    .B(_7685_),
    .Y(_7686_)
);

FILL FILL_0__18497_ (
);

AND2X2 _18362_ (
    .A(_6255__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_7273_)
);

FILL FILL412680x237120 (
);

OR2X2 _10869_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_1251_)
);

OR2X2 _10449_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_1031_)
);

OR2X2 _10029_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_811_)
);

FILL FILL_1__12952_ (
);

FILL FILL108680x79040 (
);

OR2X2 _11810_ (
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .Y(_1783_)
);

FILL FILL_0__11105_ (
);

INVX1 _19147_ (
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_8046_)
);

OR2X2 _14282_ (
    .A(vdd),
    .B(ALUOut[14]),
    .Y(_3634_)
);

FILL FILL234840x34580 (
);

FILL FILL_1__13317_ (
);

FILL FILL409640x44460 (
);

FILL FILL83600x74100 (
);

AND2X2 _15487_ (
    .A(_4154__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_4441_)
);

NAND2X1 _15067_ (
    .A(_4054_),
    .B(_4049_),
    .Y(_4055_)
);

FILL FILL_1__17990_ (
);

FILL FILL446880x256880 (
);

FILL FILL486400x365560 (
);

FILL FILL_0__16983_ (
);

FILL FILL_0__16563_ (
);

FILL FILL_0__16143_ (
);

FILL FILL378480x138320 (
);

FILL FILL_1__9700_ (
);

OR2X2 _8770_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .B(_200__bF$buf1),
    .Y(_172_)
);

FILL FILL_1__13070_ (
);

FILL FILL_0__17768_ (
);

FILL FILL231040x330980 (
);

OR2X2 _17633_ (
    .A(_6554_),
    .B(_6551_),
    .Y(_6555_)
);

FILL FILL_0__17348_ (
);

FILL FILL294880x167960 (
);

OR2X2 _17213_ (
    .A(_6138_),
    .B(_6139_),
    .Y(_6140_)
);

FILL FILL222680x207480 (
);

FILL FILL165680x19760 (
);

DFFSR _9975_ (
    .CLK(clk_bF$buf10),
    .D(_729_[3]),
    .Q(\datapath_1.regfile_1.regOut[12] [3]),
    .R(rst_bF$buf16),
    .S(vdd)
);

OR2X2 _9555_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_575_)
);

OR2X2 _9135_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_355_)
);

FILL FILL_0__8810_ (
);

FILL FILL165680x158080 (
);

FILL FILL_1__14275_ (
);

OR2X2 _18838_ (
    .A(_7710_),
    .B(_7741_),
    .Y(_7742_)
);

FILL FILL_0_BUFX2_insert550 (
);

OR2X2 _18418_ (
    .A(_7326_),
    .B(_7327_),
    .Y(_7328_)
);

FILL FILL_0_BUFX2_insert551 (
);

FILL FILL_0_BUFX2_insert552 (
);

OR2X2 _13973_ (
    .A(_3396_),
    .B(_3393_),
    .Y(\datapath_1.alu_1.ALUInB [7])
);

FILL FILL_0_BUFX2_insert554 (
);

FILL FILL_0__13268_ (
);

OR2X2 _13553_ (
    .A(ALUOut[21]),
    .B(_3079__bF$buf4),
    .Y(_3057_)
);

XOR2X1 _13133_ (
    .A(_2277_),
    .B(_2667_),
    .Y(_2685_)
);

FILL FILL_0_BUFX2_insert556 (
);

FILL FILL_0_BUFX2_insert558 (
);

AND2X2 _14758_ (
    .A(_3871_),
    .B(_3934_),
    .Y(_3870_[0])
);

DFFSR _14338_ (
    .CLK(clk_bF$buf77),
    .D(_3606_[2]),
    .Q(ALUOut[2]),
    .R(rst_bF$buf63),
    .S(vdd)
);

FILL FILL_1__16841_ (
);

FILL FILL60800x266760 (
);

FILL FILL106400x202540 (
);

FILL FILL_0__15414_ (
);

AND2X2 _18591_ (
    .A(_6262__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_7498_)
);

AND2X2 _18171_ (
    .A(_6321__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_7085_)
);

FILL FILL216600x79040 (
);

FILL FILL169480x266760 (
);

FILL FILL256880x271700 (
);

OR2X2 _10678_ (
    .A(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .B(_1190__bF$buf0),
    .Y(_1144_)
);

DFFSR _10258_ (
    .CLK(clk_bF$buf72),
    .D(_861_[28]),
    .Q(\datapath_1.regfile_1.regOut[14] [28]),
    .R(rst_bF$buf32),
    .S(vdd)
);

FILL FILL_1__17206_ (
);

FILL FILL_0__16619_ (
);

OR2X2 _16904_ (
    .A(_5835_),
    .B(_5832_),
    .Y(_5836_)
);

FILL FILL114760x316160 (
);

FILL FILL_0__11754_ (
);

FILL FILL152000x4940 (
);

AND2X2 _19376_ (
    .A(_6293__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_8271_)
);

OR2X2 _14091_ (
    .A(_3497_),
    .B(_3496_),
    .Y(_3498_)
);

DFFSR _8826_ (
    .CLK(clk_bF$buf90),
    .D(_135_[15]),
    .Q(\datapath_1.regfile_1.regOut[3] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

BUFX2 _8406_ (
    .A(_1_[14]),
    .Y(memoryAddress[14])
);

FILL FILL350360x133380 (
);

OR2X2 _12824_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2389_)
);

AND2X2 _12404_ (
    .A(_2034_),
    .B(_2033_),
    .Y(_1983_[25])
);

FILL FILL_0__12119_ (
);

FILL FILL50160x143260 (
);

FILL FILL341240x108680 (
);

OR2X2 _15296_ (
    .A(_4252_),
    .B(_4251_),
    .Y(_4253_)
);

FILL FILL_0__13900_ (
);

FILL FILL172520x103740 (
);

FILL FILL_0__16792_ (
);

FILL FILL_0__16372_ (
);

FILL FILL32680x316160 (
);

AND2X2 _13609_ (
    .A(_3089__bF$buf3),
    .B(gnd),
    .Y(_3102_)
);

FILL FILL22040x276640 (
);

FILL FILL345040x350740 (
);

FILL FILL341240x44460 (
);

FILL FILL240160x172900 (
);

FILL FILL_1__18164_ (
);

FILL FILL_0__17997_ (
);

OR2X2 _17862_ (
    .A(_6765_),
    .B(_6780_),
    .Y(_6781_)
);

AND2X2 _17442_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_6367_)
);

FILL FILL_0__17157_ (
);

AND2X2 _17022_ (
    .A(_4239__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_5952_)
);

FILL FILL_0__12292_ (
);

OR2X2 _9784_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .B(_728__bF$buf3),
    .Y(_688_)
);

OR2X2 _9364_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .B(_530__bF$buf4),
    .Y(_468_)
);

FILL FILL222680x345800 (
);

FILL FILL193800x34580 (
);

AND2X2 _18647_ (
    .A(_6328__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_7553_)
);

OR2X2 _18227_ (
    .A(_7139_),
    .B(_7136_),
    .Y(_7140_)
);

FILL FILL_0__13497_ (
);

OR2X2 _13782_ (
    .A(_3248_),
    .B(_3249_),
    .Y(_3250_)
);

FILL FILL_0__13077_ (
);

AND2X2 _13362_ (
    .A(_2900_),
    .B(_2899_),
    .Y(_2901_)
);

FILL FILL_0__19303_ (
);

FILL FILL_1__12817_ (
);

FILL FILL345040x44460 (
);

FILL FILL_0__9824_ (
);

FILL FILL_0__9404_ (
);

DFFSR _14987_ (
    .CLK(clk_bF$buf62),
    .D(_3936_[6]),
    .Q(\datapath_1.mux_iord.din0 [6]),
    .R(rst_bF$buf18),
    .S(vdd)
);

OR2X2 _14567_ (
    .A(IRWrite_bF$buf1),
    .B(\datapath_1.PCJump [25]),
    .Y(_3784_)
);

OR2X2 _14147_ (
    .A(\datapath_1.Data [1]),
    .B(_3605__bF$buf1),
    .Y(_3543_)
);

FILL FILL231800x49400 (
);

FILL FILL_0__15643_ (
);

FILL FILL250800x227240 (
);

FILL FILL46360x49400 (
);

FILL FILL197600x34580 (
);

AND2X2 _10487_ (
    .A(_1056_),
    .B(_1055_),
    .Y(_993_[31])
);

AND2X2 _10067_ (
    .A(_836_),
    .B(_835_),
    .Y(_795_[20])
);

FILL FILL_1__12150_ (
);

FILL FILL_0__16848_ (
);

OR2X2 _16713_ (
    .A(_5647_),
    .B(_5640_),
    .Y(_5648_)
);

FILL FILL_0__16008_ (
);

FILL FILL_0__11983_ (
);

FILL FILL_0__11563_ (
);

OR2X2 _19185_ (
    .A(_8079_),
    .B(_8082_),
    .Y(_8083_)
);

FILL FILL368600x217360 (
);

OR2X2 _8635_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .B(_134__bF$buf3),
    .Y(_102_)
);

FILL FILL31920x167960 (
);

FILL FILL303240x74100 (
);

OR2X2 _17918_ (
    .A(_6832_),
    .B(_6835_),
    .Y(_6836_)
);

FILL FILL_0__12768_ (
);

OR2X2 _12633_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(_2197_),
    .Y(_2198_)
);

OR2X2 _12213_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_1927_)
);

OR2X2 _13838_ (
    .A(\datapath_1.a [7]),
    .B(_3342__bF$buf2),
    .Y(_3292_)
);

NAND2X1 _13418_ (
    .A(_2388_),
    .B(_2379__bF$buf2),
    .Y(_2953_)
);

FILL FILL132240x64220 (
);

FILL FILL_0__14914_ (
);

FILL FILL_0__17386_ (
);

AND2X2 _17671_ (
    .A(_6206__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_6592_)
);

OR2X2 _17251_ (
    .A(_6176_),
    .B(_6177_),
    .Y(_6178_)
);

FILL FILL294120x335920 (
);

FILL FILL129200x247000 (
);

DFFSR _9593_ (
    .CLK(clk_bF$buf22),
    .D(_531_[8]),
    .Q(\datapath_1.regfile_1.regOut[9] [8]),
    .R(rst_bF$buf74),
    .S(vdd)
);

FILL FILL_1__16706_ (
);

AND2X2 _9173_ (
    .A(_380_),
    .B(_379_),
    .Y(_333_[23])
);

FILL FILL_1__11841_ (
);

FILL FILL_1__19178_ (
);

FILL FILL_0__10834_ (
);

FILL FILL229520x340860 (
);

OR2X2 _18876_ (
    .A(_7778_),
    .B(_7777_),
    .Y(_7779_)
);

FILL FILL_0_BUFX2_insert930 (
);

FILL FILL_0_BUFX2_insert931 (
);

OR2X2 _18456_ (
    .A(_7363_),
    .B(_7364_),
    .Y(_7365_)
);

AND2X2 _18036_ (
    .A(_6300__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_6952_)
);

FILL FILL_0_BUFX2_insert933 (
);

OR2X2 _13591_ (
    .A(_3082_),
    .B(_3085_),
    .Y(_3086_)
);

FILL FILL_0_BUFX2_insert935 (
);

INVX1 _13171_ (
    .A(_2717_),
    .Y(_2721_)
);

FILL FILL_0_BUFX2_insert937 (
);

FILL FILL447640x143260 (
);

FILL FILL_0_BUFX2_insert939 (
);

FILL FILL_0__19112_ (
);

FILL FILL430160x227240 (
);

FILL FILL367080x0 (
);

FILL FILL_1__12206_ (
);

FILL FILL474240x83980 (
);

FILL FILL_0__9633_ (
);

OR2X2 _11904_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_1781_)
);

FILL FILL270560x49400 (
);

FILL FILL333640x261820 (
);

OR2X2 _14796_ (
    .A(\datapath_1.rd2 [13]),
    .B(_3935__bF$buf1),
    .Y(_3897_)
);

OR2X2 _14376_ (
    .A(memoryOutData[2]),
    .B(_3737__bF$buf3),
    .Y(_3677_)
);

FILL FILL47120x247000 (
);

FILL FILL_0__15452_ (
);

FILL FILL_0__15032_ (
);

FILL FILL_1__17664_ (
);

OR2X2 _10296_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_949_)
);

FILL FILL_0__16657_ (
);

OR2X2 _16942_ (
    .A(_5873_),
    .B(_5872_),
    .Y(_5874_)
);

AND2X2 _16522_ (
    .A(_4203__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_5460_)
);

FILL FILL_0__16237_ (
);

OR2X2 _16102_ (
    .A(_5045_),
    .B(_5046_),
    .Y(_5047_)
);

FILL FILL_0__11372_ (
);

AND2X2 _8864_ (
    .A(_214_),
    .B(_213_),
    .Y(_201_[6])
);

BUFX2 _8444_ (
    .A(_2_[20]),
    .Y(memoryWriteData[20])
);

FILL FILL_1__18029_ (
);

AND2X2 _17727_ (
    .A(_6323__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_6648_)
);

AND2X2 _17307_ (
    .A(_6232__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [0]),
    .Y(_6233_)
);

FILL FILL_0__12997_ (
);

OR2X2 _12862_ (
    .A(_2221_),
    .B(_2222_),
    .Y(_2427_)
);

DFFSR _12442_ (
    .CLK(clk_bF$buf69),
    .D(_1983_[19]),
    .Q(\datapath_1.regfile_1.regOut[31] [19]),
    .R(rst_bF$buf79),
    .S(vdd)
);

FILL FILL_0__12157_ (
);

OR2X2 _12022_ (
    .A(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .B(_1850__bF$buf2),
    .Y(_1840_)
);

FILL FILL_0__18803_ (
);

OR2X2 _9649_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .B(_662__bF$buf4),
    .Y(_618_)
);

DFFSR _9229_ (
    .CLK(clk_bF$buf56),
    .D(_333_[31]),
    .Q(\datapath_1.regfile_1.regOut[6] [31]),
    .R(rst_bF$buf30),
    .S(vdd)
);

FILL FILL323760x59280 (
);

FILL FILL_0__8904_ (
);

AND2X2 _13647_ (
    .A(_3081__bF$buf0),
    .B(ALUOut[8]),
    .Y(_3134_)
);

AND2X2 _13227_ (
    .A(_2773_),
    .B(_2248_),
    .Y(_2774_)
);

FILL FILL_1__15310_ (
);

FILL FILL_0__14303_ (
);

AND2X2 _17480_ (
    .A(_6232__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .Y(_6404_)
);

AND2X2 _17060_ (
    .A(_4236__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_5990_)
);

FILL FILL34960x44460 (
);

FILL FILL_0_CLKBUF1_insert160 (
);

FILL FILL_1__11230_ (
);

FILL FILL_0_CLKBUF1_insert162 (
);

FILL FILL_0__15928_ (
);

FILL FILL_0__15508_ (
);

FILL FILL_0_CLKBUF1_insert164 (
);

FILL FILL_0_CLKBUF1_insert166 (
);

FILL FILL_0_CLKBUF1_insert168 (
);

FILL FILL_0_CLKBUF1_insert169 (
);

AND2X2 _18685_ (
    .A(_6326__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_7591_)
);

OR2X2 _18265_ (
    .A(_7175_),
    .B(_7176_),
    .Y(_7177_)
);

FILL FILL379240x118560 (
);

FILL FILL466640x123500 (
);

FILL FILL202160x301340 (
);

FILL FILL171000x49400 (
);

FILL FILL_0__11848_ (
);

FILL FILL_0__9442_ (
);

FILL FILL_0__11428_ (
);

FILL FILL_0__9022_ (
);

OR2X2 _11713_ (
    .A(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .B(_1718__bF$buf1),
    .Y(_1674_)
);

OR2X2 _14185_ (
    .A(MemToReg_bF$buf2),
    .B(ALUOut[14]),
    .Y(_3568_)
);

FILL FILL200640x44460 (
);

FILL FILL439280x34580 (
);

FILL FILL_0__15681_ (
);

FILL FILL_0__15261_ (
);

FILL FILL483360x360620 (
);

FILL FILL_1_BUFX2_insert480 (
);

AOI21X1 _12918_ (
    .A(_2481_),
    .B(_2478_),
    .C(_2482_),
    .Y(_2483_)
);

FILL FILL_1_BUFX2_insert482 (
);

FILL FILL367080x98800 (
);

FILL FILL_1_BUFX2_insert484 (
);

FILL FILL266000x74100 (
);

FILL FILL_0__16886_ (
);

OR2X2 _16751_ (
    .A(_5685_),
    .B(_5682_),
    .Y(_5686_)
);

FILL FILL_0__16466_ (
);

AND2X2 _16331_ (
    .A(_4239__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_5272_)
);

FILL FILL_0__11181_ (
);

OR2X2 _8673_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_127_)
);

FILL FILL50160x306280 (
);

FILL FILL_1__10921_ (
);

FILL FILL_1__18678_ (
);

FILL FILL_1__13393_ (
);

OR2X2 _17956_ (
    .A(_6872_),
    .B(_6871_),
    .Y(_6873_)
);

OR2X2 _17536_ (
    .A(_6459_),
    .B(_6452_),
    .Y(_6460_)
);

FILL FILL234840x167960 (
);

OR2X2 _17116_ (
    .A(_6043_),
    .B(_6044_),
    .Y(_6045_)
);

INVX1 _12671_ (
    .A(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2236_)
);

AND2X2 _12251_ (
    .A(_1952_),
    .B(_1951_),
    .Y(_1917_[17])
);

FILL FILL367080x163020 (
);

FILL FILL_0__18612_ (
);

FILL FILL371640x227240 (
);

AND2X2 _9878_ (
    .A(_730_),
    .B(_793_),
    .Y(_729_[0])
);

DFFSR _9458_ (
    .CLK(clk_bF$buf17),
    .D(_465_[2]),
    .Q(\datapath_1.regfile_1.regOut[8] [2]),
    .R(rst_bF$buf113),
    .S(vdd)
);

AND2X2 _9038_ (
    .A(_310_),
    .B(_309_),
    .Y(_267_[21])
);

FILL FILL272080x123500 (
);

OR2X2 _13876_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.mux_iord.din0 [20]),
    .Y(_3317_)
);

AND2X2 _13456_ (
    .A(_2988_),
    .B(_2935_),
    .Y(_2989_)
);

FILL FILL211280x232180 (
);

AOI22X1 _13036_ (
    .A(_2592_),
    .B(_2379__bF$buf0),
    .C(_2593_),
    .D(_2334_),
    .Y(_2594_)
);

FILL FILL_0__14952_ (
);

FILL FILL_0__14112_ (
);

FILL FILL183160x286520 (
);

FILL FILL_0__9918_ (
);

FILL FILL93480x59280 (
);

FILL FILL_1__10098_ (
);

FILL FILL158840x29640 (
);

FILL FILL_0__15737_ (
);

FILL FILL505400x291460 (
);

FILL FILL_0__15317_ (
);

OR2X2 _15602_ (
    .A(_4554_),
    .B(_4553_),
    .Y(_4555_)
);

FILL FILL_0__10872_ (
);

FILL FILL_0__10452_ (
);

OR2X2 _18494_ (
    .A(_7401_),
    .B(_7402_),
    .Y(_7403_)
);

OR2X2 _18074_ (
    .A(_6988_),
    .B(_6987_),
    .Y(_6989_)
);

FILL FILL_0__19150_ (
);

FILL FILL75240x345800 (
);

FILL FILL_1__17529_ (
);

FILL FILL180120x182780 (
);

FILL FILL53960x14820 (
);

FILL FILL212040x9880 (
);

OR2X2 _16807_ (
    .A(_5737_),
    .B(_5740_),
    .Y(_5741_)
);

FILL FILL126920x276640 (
);

FILL FILL_0__9671_ (
);

AND2X2 _11942_ (
    .A(_1786_),
    .B(_1849_),
    .Y(_1785_[0])
);

FILL FILL_0__9251_ (
);

FILL FILL282720x59280 (
);

FILL FILL_0__11237_ (
);

DFFSR _11522_ (
    .CLK(clk_bF$buf51),
    .D(_1521_[2]),
    .Q(\datapath_1.regfile_1.regOut[24] [2]),
    .R(rst_bF$buf12),
    .S(vdd)
);

AND2X2 _11102_ (
    .A(_1366_),
    .B(_1365_),
    .Y(_1323_[21])
);

OR2X2 _19279_ (
    .A(_8174_),
    .B(_8175_),
    .Y(_8176_)
);

AND2X2 _8729_ (
    .A(_144_),
    .B(_143_),
    .Y(_135_[4])
);

FILL FILL433960x103740 (
);

FILL FILL457520x69160 (
);

FILL FILL_0__15490_ (
);

FILL FILL_0__15070_ (
);

FILL FILL_1__13869_ (
);

INVX1 _12727_ (
    .A(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2292_)
);

DFFSR _12307_ (
    .CLK(clk_bF$buf85),
    .D(_1917_[13]),
    .Q(\datapath_1.regfile_1.regOut[30] [13]),
    .R(rst_bF$buf60),
    .S(vdd)
);

FILL FILL410400x39520 (
);

AND2X2 _15199_ (
    .A(_4133_),
    .B(_4139_),
    .Y(_4157_)
);

FILL FILL_0__13803_ (
);

FILL FILL_1__17282_ (
);

AND2X2 _16980_ (
    .A(_4214__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_5911_)
);

AND2X2 _16560_ (
    .A(_4142__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_5498_)
);

OR2X2 _16140_ (
    .A(_5083_),
    .B(_5082_),
    .Y(_5084_)
);

FILL FILL_1__9832_ (
);

FILL FILL473480x103740 (
);

OR2X2 _8482_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .B(_68__bF$buf1),
    .Y(_20_)
);

FILL FILL123120x54340 (
);

FILL FILL367080x256880 (
);

FILL FILL505400x64220 (
);

OR2X2 _17765_ (
    .A(_6684_),
    .B(_6671_),
    .Y(_6685_)
);

AND2X2 _17345_ (
    .A(_6270_),
    .B(_6201_),
    .Y(_6271_)
);

AND2X2 _12480_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2072_)
);

DFFSR _12060_ (
    .CLK(clk_bF$buf35),
    .D(_1785_[24]),
    .Q(\datapath_1.regfile_1.regOut[28] [24]),
    .R(rst_bF$buf6),
    .S(vdd)
);

FILL FILL110200x177840 (
);

FILL FILL_0__18841_ (
);

FILL FILL_0__18421_ (
);

FILL FILL_0__18001_ (
);

OR2X2 _9687_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_643_)
);

OR2X2 _9267_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_423_)
);

FILL FILL_1_CLKBUF1_insert190 (
);

FILL FILL_1_CLKBUF1_insert198 (
);

FILL FILL_0__8522_ (
);

FILL FILL_0__10928_ (
);

FILL FILL272840x4940 (
);

AND2X2 _13685_ (
    .A(_3087__bF$buf3),
    .B(\datapath_1.ALUResult [13]),
    .Y(_3167_)
);

OR2X2 _13265_ (
    .A(_2157__bF$buf3),
    .B(_2808_),
    .Y(_2809_)
);

FILL FILL_0__14761_ (
);

FILL FILL_0__9307_ (
);

FILL FILL291840x4940 (
);

FILL FILL173280x163020 (
);

FILL FILL447640x306280 (
);

FILL FILL_1__16133_ (
);

FILL FILL351120x251940 (
);

FILL FILL25080x128440 (
);

FILL FILL_0__15966_ (
);

OR2X2 _15831_ (
    .A(_4776_),
    .B(_4779_),
    .Y(_4780_)
);

FILL FILL_0__15126_ (
);

AND2X2 _15411_ (
    .A(_4214__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_4367_)
);

FILL FILL_0__10681_ (
);

FILL FILL433960x330980 (
);

FILL FILL61560x301340 (
);

FILL FILL281200x256880 (
);

FILL FILL42560x138320 (
);

FILL FILL365560x212420 (
);

FILL FILL_1__17758_ (
);

OR2X2 _16616_ (
    .A(_5552_),
    .B(_5545_),
    .Y(_5553_)
);

FILL FILL295640x217360 (
);

FILL FILL_0__11886_ (
);

OR2X2 _11751_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_1699_)
);

FILL FILL_0__9060_ (
);

FILL FILL_0__11046_ (
);

OR2X2 _11331_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_1479_)
);

OR2X2 _19088_ (
    .A(_7987_),
    .B(_7984_),
    .Y(_7988_)
);

FILL FILL276640x375440 (
);

DFFSR _8958_ (
    .CLK(clk_bF$buf91),
    .D(_201_[18]),
    .Q(\datapath_1.regfile_1.regOut[4] [18]),
    .R(rst_bF$buf50),
    .S(vdd)
);

OR2X2 _8538_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_57_)
);

FILL FILL265240x39520 (
);

FILL FILL181640x335920 (
);

FILL FILL_1__13258_ (
);

FILL FILL_1_BUFX2_insert860 (
);

AOI21X1 _12956_ (
    .A(ALUControl[1]),
    .B(_2353_),
    .C(_2518_),
    .Y(_2519_)
);

FILL FILL_1_BUFX2_insert862 (
);

FILL FILL392920x54340 (
);

OR2X2 _12536_ (
    .A(IRWrite_bF$buf2),
    .B(_2125_),
    .Y(_2126_)
);

FILL FILL_1_BUFX2_insert864 (
);

AND2X2 _12116_ (
    .A(_1882_),
    .B(_1881_),
    .Y(_1851_[15])
);

FILL FILL_0__16084_ (
);

FILL FILL_1__9641_ (
);

FILL FILL_1__15824_ (
);

FILL FILL_0__14817_ (
);

BUFX2 BUFX2_insert530 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf109)
);

BUFX2 BUFX2_insert531 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf108)
);

BUFX2 BUFX2_insert532 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf107)
);

BUFX2 BUFX2_insert533 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf106)
);

BUFX2 BUFX2_insert534 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf105)
);

OR2X2 _17994_ (
    .A(_6876_),
    .B(_6910_),
    .Y(_6911_)
);

AND2X2 _17574_ (
    .A(_6229__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_6497_)
);

BUFX2 BUFX2_insert535 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf104)
);

FILL FILL_0__17289_ (
);

BUFX2 BUFX2_insert536 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf103)
);

AND2X2 _17154_ (
    .A(_4151__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_6082_)
);

BUFX2 BUFX2_insert537 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf102)
);

BUFX2 BUFX2_insert538 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf101)
);

BUFX2 BUFX2_insert539 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf100)
);

FILL FILL321480x148200 (
);

FILL FILL_0__18650_ (
);

FILL FILL_0__18230_ (
);

OR2X2 _9496_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .B(_596__bF$buf3),
    .Y(_536_)
);

DFFSR _9076_ (
    .CLK(clk_bF$buf66),
    .D(_267_[7]),
    .Q(\datapath_1.regfile_1.regOut[5] [7]),
    .R(rst_bF$buf69),
    .S(vdd)
);

FILL FILL_0__8751_ (
);

OR2X2 _10602_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_1113_)
);

FILL FILL_0_BUFX2_insert50 (
);

AND2X2 _18779_ (
    .A(_6271__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_7683_)
);

FILL FILL_0_BUFX2_insert52 (
);

AND2X2 _18359_ (
    .A(_6221__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_7270_)
);

FILL FILL_0_BUFX2_insert54 (
);

FILL FILL_0_BUFX2_insert56 (
);

AND2X2 _13494_ (
    .A(_3017_),
    .B(_3016_),
    .Y(_1_[1])
);

NOR3X1 _13074_ (
    .A(_2629_),
    .B(_2626_),
    .C(_2627_),
    .Y(_2630_)
);

FILL FILL_0_BUFX2_insert58 (
);

FILL FILL_0_BUFX2_insert59 (
);

FILL FILL_0__19015_ (
);

NOR2X1 _19300_ (
    .A(_6310__bF$buf4),
    .B(_8195_),
    .Y(_8196_)
);

FILL FILL57760x103740 (
);

FILL FILL_0__14150_ (
);

FILL FILL_1__12529_ (
);

FILL FILL_0__9956_ (
);

FILL FILL_0__9536_ (
);

FILL FILL_0__9116_ (
);

DFFSR _11807_ (
    .CLK(clk_bF$buf11),
    .D(_1653_[29]),
    .Q(\datapath_1.regfile_1.regOut[26] [29]),
    .R(rst_bF$buf111),
    .S(vdd)
);

FILL FILL69920x247000 (
);

OR2X2 _14699_ (
    .A(vdd),
    .B(\datapath_1.a [24]),
    .Y(_3852_)
);

OR2X2 _14279_ (
    .A(vdd),
    .B(ALUOut[13]),
    .Y(_3632_)
);

FILL FILL_1__16782_ (
);

FILL FILL_0__15775_ (
);

FILL FILL_0__15355_ (
);

OR2X2 _15640_ (
    .A(_4591_),
    .B(_4584_),
    .Y(_4592_)
);

AND2X2 _15220_ (
    .A(_4177__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_4178_)
);

FILL FILL410400x321100 (
);

FILL FILL74480x340860 (
);

FILL FILL_0__10070_ (
);

FILL FILL_1__8912_ (
);

AND2X2 _10199_ (
    .A(_904_),
    .B(_903_),
    .Y(_861_[21])
);

FILL FILL_1__17147_ (
);

FILL FILL_1__12282_ (
);

AND2X2 _16845_ (
    .A(_4214__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_5778_)
);

AND2X2 _16425_ (
    .A(_4214__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_5365_)
);

AND2X2 _16005_ (
    .A(_4172__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_4951_)
);

OR2X2 _11980_ (
    .A(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .B(_1850__bF$buf4),
    .Y(_1812_)
);

FILL FILL_0__11695_ (
);

OR2X2 _11560_ (
    .A(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .B(_1652__bF$buf1),
    .Y(_1592_)
);

DFFSR _11140_ (
    .CLK(clk_bF$buf48),
    .D(_1323_[7]),
    .Q(\datapath_1.regfile_1.regOut[21] [7]),
    .R(rst_bF$buf48),
    .S(vdd)
);

FILL FILL252320x291460 (
);

FILL FILL496280x148200 (
);

FILL FILL_0__17921_ (
);

OR2X2 _8767_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .B(_200__bF$buf0),
    .Y(_170_)
);

FILL FILL418760x207480 (
);

FILL FILL_1__13487_ (
);

OR2X2 _12765_ (
    .A(_2329_),
    .B(_2328_),
    .Y(_2330_)
);

OR2X2 _12345_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_1995_)
);

FILL FILL135280x360620 (
);

FILL FILL425600x177840 (
);

FILL FILL_0__13421_ (
);

FILL FILL_0__13001_ (
);

FILL FILL321480x375440 (
);

FILL FILL_0__8807_ (
);

FILL FILL_1__9030_ (
);

FILL FILL_0__14626_ (
);

AND2X2 _14911_ (
    .A(_3953_),
    .B(_3952_),
    .Y(_3936_[8])
);

FILL FILL_0__14206_ (
);

OR2X2 _17383_ (
    .A(_6308_),
    .B(_6257_),
    .Y(_6309_)
);

FILL FILL_0__17098_ (
);

FILL FILL9120x167960 (
);

FILL FILL333640x19760 (
);

FILL FILL_1__11973_ (
);

FILL FILL_0__10966_ (
);

OR2X2 _10831_ (
    .A(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .B(_1256__bF$buf2),
    .Y(_1226_)
);

OR2X2 _10411_ (
    .A(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .B(_1058__bF$buf4),
    .Y(_1006_)
);

AND2X2 _18588_ (
    .A(_6247__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_7495_)
);

OR2X2 _18168_ (
    .A(_7080_),
    .B(_7081_),
    .Y(_7082_)
);

FILL FILL_0__19244_ (
);

FILL FILL253840x34580 (
);

FILL FILL_1__12338_ (
);

FILL FILL_0__9765_ (
);

OR2X2 _11616_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_1629_)
);

FILL FILL381520x232180 (
);

FILL FILL428640x44460 (
);

OR2X2 _14088_ (
    .A(_3493_),
    .B(_3494_),
    .Y(_3495_)
);

FILL FILL_0__15584_ (
);

FILL FILL414960x237120 (
);

FILL FILL_1__8721_ (
);

FILL FILL404320x197600 (
);

FILL FILL24320x69160 (
);

FILL FILL_1__17796_ (
);

FILL FILL285000x247000 (
);

FILL FILL_1__12091_ (
);

AND2X2 _16654_ (
    .A(_4154__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_5590_)
);

FILL FILL_0__16369_ (
);

AND2X2 _16234_ (
    .A(_4239__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_5177_)
);

FILL FILL281960x311220 (
);

FILL FILL440040x276640 (
);

FILL FILL_1__9926_ (
);

FILL FILL_0__17730_ (
);

FILL FILL_0__17310_ (
);

FILL FILL268280x222300 (
);

AND2X2 _8996_ (
    .A(_282_),
    .B(_281_),
    .Y(_267_[7])
);

DFFSR _8576_ (
    .CLK(clk_bF$buf84),
    .D(_3_[23]),
    .Q(\datapath_1.regfile_1.regOut[1] [23]),
    .R(rst_bF$buf47),
    .S(vdd)
);

FILL FILL167960x69160 (
);

FILL FILL279680x291460 (
);

OR2X2 _17859_ (
    .A(_6777_),
    .B(_6776_),
    .Y(_6778_)
);

OR2X2 _17439_ (
    .A(_6363_),
    .B(_6356_),
    .Y(_6364_)
);

AND2X2 _17019_ (
    .A(_4217__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_5949_)
);

OR2X2 _12994_ (
    .A(_2554_),
    .B(_2475_),
    .Y(_2555_)
);

FILL FILL_0__12289_ (
);

AND2X2 _12574_ (
    .A(_2146_),
    .B(_2144_),
    .Y(_2143_[0])
);

OR2X2 _12154_ (
    .A(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .B(_1916__bF$buf3),
    .Y(_1908_)
);

FILL FILL_0__18935_ (
);

NOR2X1 _18800_ (
    .A(_6310__bF$buf1),
    .B(_7703_),
    .Y(_7704_)
);

FILL FILL_0__18515_ (
);

FILL FILL66120x187720 (
);

FILL FILL_0__13650_ (
);

FILL FILL_0__13230_ (
);

FILL FILL_1__11609_ (
);

OR2X2 _13779_ (
    .A(_3247_),
    .B(_3244_),
    .Y(\datapath_1.mux_pcsrc.dout [26])
);

AOI21X1 _13359_ (
    .A(_2896_),
    .B(_2897_),
    .C(_2895_),
    .Y(_2898_)
);

OR2X2 _14720_ (
    .A(vdd),
    .B(\datapath_1.a [31]),
    .Y(_3866_)
);

FILL FILL_0__14435_ (
);

OR2X2 _14300_ (
    .A(vdd),
    .B(ALUOut[20]),
    .Y(_3646_)
);

BUFX2 BUFX2_insert910 (
    .A(_6293_),
    .Y(_6293__bF$buf2)
);

BUFX2 BUFX2_insert911 (
    .A(_6293_),
    .Y(_6293__bF$buf1)
);

BUFX2 BUFX2_insert912 (
    .A(_6293_),
    .Y(_6293__bF$buf0)
);

BUFX2 BUFX2_insert913 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf4 )
);

BUFX2 BUFX2_insert914 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf3 )
);

BUFX2 BUFX2_insert915 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf2 )
);

OR2X2 _17192_ (
    .A(_6119_),
    .B(_6112_),
    .Y(_6120_)
);

BUFX2 BUFX2_insert916 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf1 )
);

BUFX2 BUFX2_insert917 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf0 )
);

BUFX2 BUFX2_insert918 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf4 )
);

BUFX2 BUFX2_insert919 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf3 )
);

FILL FILL176320x281580 (
);

FILL FILL_1__16647_ (
);

FILL FILL_1__16227_ (
);

FILL FILL_1__11362_ (
);

OR2X2 _15925_ (
    .A(_4871_),
    .B(_4872_),
    .Y(_4873_)
);

AND2X2 _15505_ (
    .A(_4151__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_4459_)
);

DFFSR _10640_ (
    .CLK(clk_bF$buf26),
    .D(_1059_[23]),
    .Q(\datapath_1.regfile_1.regOut[17] [23]),
    .R(rst_bF$buf94),
    .S(vdd)
);

AND2X2 _10220_ (
    .A(_918_),
    .B(_917_),
    .Y(_861_[28])
);

FILL FILL212040x79040 (
);

AND2X2 _18397_ (
    .A(_6211__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_7307_)
);

FILL FILL358720x192660 (
);

FILL FILL173280x326040 (
);

FILL FILL_0__19053_ (
);

FILL FILL_1__12987_ (
);

FILL FILL_0__9574_ (
);

OR2X2 _11845_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .B(_1784__bF$buf4),
    .Y(_1742_)
);

FILL FILL_0__9154_ (
);

FILL FILL86640x69160 (
);

OR2X2 _11425_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(_1586__bF$buf4),
    .Y(_1522_)
);

DFFSR _11005_ (
    .CLK(clk_bF$buf47),
    .D(_1257_[1]),
    .Q(\datapath_1.regfile_1.regOut[20] [1]),
    .R(rst_bF$buf103),
    .S(vdd)
);

FILL FILL_0__12921_ (
);

FILL FILL_0__12501_ (
);

FILL FILL423320x79040 (
);

FILL FILL440040x29640 (
);

FILL FILL146680x49400 (
);

FILL FILL_1__8530_ (
);

FILL FILL372400x345800 (
);

FILL FILL_0__16598_ (
);

AND2X2 _16883_ (
    .A(_4230__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_5816_)
);

FILL FILL_0__16178_ (
);

OR2X2 _16463_ (
    .A(_5401_),
    .B(_5400_),
    .Y(_5402_)
);

OR2X2 _16043_ (
    .A(_4988_),
    .B(_4987_),
    .Y(_4989_)
);

FILL FILL213560x88920 (
);

FILL FILL203680x227240 (
);

FILL FILL467400x29640 (
);

OR2X2 _17668_ (
    .A(_6558_),
    .B(_6589_),
    .Y(_6590_)
);

FILL FILL343520x108680 (
);

OR2X2 _17248_ (
    .A(_6174_),
    .B(_6171_),
    .Y(_6175_)
);

FILL FILL430920x113620 (
);

AND2X2 _12383_ (
    .A(_2020_),
    .B(_2019_),
    .Y(_1983_[18])
);

FILL FILL_0__12098_ (
);

FILL FILL174800x103740 (
);

FILL FILL_0__18744_ (
);

FILL FILL408880x222300 (
);

FILL FILL430160x340860 (
);

FILL FILL_0__8845_ (
);

FILL FILL347320x350740 (
);

INVX1 _13588_ (
    .A(ALUOp[0]),
    .Y(_3083_)
);

INVX1 _13168_ (
    .A(_2283_),
    .Y(_2718_)
);

FILL FILL217360x88920 (
);

FILL FILL481840x79040 (
);

FILL FILL_1__15251_ (
);

FILL FILL_0__19109_ (
);

FILL FILL_0__14244_ (
);

FILL FILL224960x345800 (
);

FILL FILL247000x83980 (
);

FILL FILL113240x163020 (
);

FILL FILL_1__16876_ (
);

FILL FILL_0__15869_ (
);

FILL FILL_0__15449_ (
);

OR2X2 _15734_ (
    .A(_4681_),
    .B(_4684_),
    .Y(_4685_)
);

AND2X2 _15314_ (
    .A(_4225__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_4271_)
);

FILL FILL_0__10584_ (
);

FILL FILL193040x34580 (
);

BUFX2 BUFX2_insert60 (
    .A(_4217_),
    .Y(_4217__bF$buf4)
);

BUFX2 BUFX2_insert61 (
    .A(_4217_),
    .Y(_4217__bF$buf3)
);

BUFX2 BUFX2_insert62 (
    .A(_4217_),
    .Y(_4217__bF$buf2)
);

FILL FILL370880x9880 (
);

BUFX2 BUFX2_insert63 (
    .A(_4217_),
    .Y(_4217__bF$buf1)
);

BUFX2 BUFX2_insert64 (
    .A(_4217_),
    .Y(_4217__bF$buf0)
);

FILL FILL_0__16810_ (
);

BUFX2 BUFX2_insert65 (
    .A(_4158_),
    .Y(_4158__bF$buf4)
);

BUFX2 BUFX2_insert66 (
    .A(_4158_),
    .Y(_4158__bF$buf3)
);

BUFX2 BUFX2_insert67 (
    .A(_4158_),
    .Y(_4158__bF$buf2)
);

BUFX2 BUFX2_insert68 (
    .A(_4158_),
    .Y(_4158__bF$buf1)
);

BUFX2 BUFX2_insert69 (
    .A(_4158_),
    .Y(_4158__bF$buf0)
);

FILL FILL_0__19282_ (
);

FILL FILL485640x79040 (
);

OR2X2 _16939_ (
    .A(_5869_),
    .B(_5870_),
    .Y(_5871_)
);

OR2X2 _16519_ (
    .A(_5455_),
    .B(_5456_),
    .Y(_5457_)
);

FILL FILL_0__9383_ (
);

DFFSR _11654_ (
    .CLK(clk_bF$buf66),
    .D(_1587_[5]),
    .Q(\datapath_1.regfile_1.regOut[25] [5]),
    .R(rst_bF$buf80),
    .S(vdd)
);

AND2X2 _11234_ (
    .A(_1434_),
    .B(_1433_),
    .Y(_1389_[22])
);

FILL FILL231040x49400 (
);

OR2X2 _9802_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .B(_728__bF$buf3),
    .Y(_700_)
);

OR2X2 _12859_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2424_)
);

DFFSR _12439_ (
    .CLK(clk_bF$buf78),
    .D(_1983_[16]),
    .Q(\datapath_1.regfile_1.regOut[31] [16]),
    .R(rst_bF$buf110),
    .S(vdd)
);

OR2X2 _12019_ (
    .A(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .B(_1850__bF$buf0),
    .Y(_1838_)
);

FILL FILL_0__13935_ (
);

FILL FILL_0__13515_ (
);

OR2X2 _13800_ (
    .A(_3265_),
    .B(_3262_),
    .Y(\datapath_1.mux_pcsrc.dout [29])
);

AND2X2 _16692_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_5628_)
);

OR2X2 _16272_ (
    .A(_5210_),
    .B(_5213_),
    .Y(_5214_)
);

FILL FILL_1__9964_ (
);

FILL FILL_1__10862_ (
);

FILL FILL258400x49400 (
);

FILL FILL_1__18199_ (
);

AND2X2 _17897_ (
    .A(_6271__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_6815_)
);

AND2X2 _17477_ (
    .A(_6216__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_6401_)
);

AND2X2 _17057_ (
    .A(_4158__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_5987_)
);

FILL FILL4560x192660 (
);

DFFSR _12192_ (
    .CLK(clk_bF$buf14),
    .D(_1851_[27]),
    .Q(\datapath_1.regfile_1.regOut[29] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

FILL FILL300200x182780 (
);

FILL FILL_0__18133_ (
);

OR2X2 _9399_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_491_)
);

FILL FILL_0__8654_ (
);

FILL FILL92720x93860 (
);

AND2X2 _10925_ (
    .A(_1268_),
    .B(_1267_),
    .Y(_1257_[5])
);

DFFSR _10505_ (
    .CLK(clk_bF$buf109),
    .D(_993_[17]),
    .Q(\datapath_1.regfile_1.regOut[16] [17]),
    .R(rst_bF$buf84),
    .S(vdd)
);

AND2X2 _13397_ (
    .A(_2933_),
    .B(_2928_),
    .Y(_2934_)
);

FILL FILL_0__19338_ (
);

AND2X2 _19203_ (
    .A(_6302__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_8101_)
);

FILL FILL_0__14893_ (
);

FILL FILL28120x316160 (
);

FILL FILL_1__16265_ (
);

AND2X2 _15963_ (
    .A(_4175__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_4910_)
);

OR2X2 _15543_ (
    .A(_4496_),
    .B(_4489_),
    .Y(_4497_)
);

AND2X2 _15123_ (
    .A(_4100_),
    .B(_4035_),
    .Y(_4101_)
);

FILL FILL_0__10393_ (
);

FILL FILL_0__19091_ (
);

FILL FILL293360x49400 (
);

FILL FILL504640x266760 (
);

AND2X2 _16748_ (
    .A(_4228__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_5683_)
);

OR2X2 _16328_ (
    .A(_5265_),
    .B(_5268_),
    .Y(_5269_)
);

OR2X2 _11883_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_1767_)
);

OR2X2 _11463_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_1547_)
);

FILL FILL_1__18411_ (
);

OR2X2 _11043_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_1327_)
);

FILL FILL_0__17404_ (
);

DFFSR _9611_ (
    .CLK(clk_bF$buf86),
    .D(_531_[26]),
    .Q(\datapath_1.regfile_1.regOut[9] [26]),
    .R(rst_bF$buf42),
    .S(vdd)
);

FILL FILL197600x148200 (
);

AND2X2 _12668_ (
    .A(_2232_),
    .B(_2228_),
    .Y(_2233_)
);

AND2X2 _12248_ (
    .A(_1950_),
    .B(_1949_),
    .Y(_1917_[16])
);

FILL FILL_0__18609_ (
);

FILL FILL_0__13744_ (
);

FILL FILL_0__13324_ (
);

FILL FILL148960x335920 (
);

AND2X2 _16081_ (
    .A(_4214__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_5026_)
);

FILL FILL407360x232180 (
);

FILL FILL_1__9773_ (
);

FILL FILL_1__15116_ (
);

FILL FILL387600x88920 (
);

FILL FILL_1__10671_ (
);

FILL FILL_0__14949_ (
);

OR2X2 _14814_ (
    .A(\datapath_1.rd2 [19]),
    .B(_3935__bF$buf4),
    .Y(_3909_)
);

FILL FILL_0__14529_ (
);

FILL FILL_0__14109_ (
);

AND2X2 _17286_ (
    .A(_6211__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_6212_)
);

FILL FILL12160x202540 (
);

FILL FILL346560x59280 (
);

FILL FILL_0__18782_ (
);

FILL FILL_0__18362_ (
);

FILL FILL_1__11036_ (
);

FILL FILL_0__8463_ (
);

FILL FILL_0__10869_ (
);

OR2X2 _10734_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_1181_)
);

FILL FILL_0__10029_ (
);

OR2X2 _10314_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_961_)
);

FILL FILL310080x266760 (
);

FILL FILL237880x316160 (
);

FILL FILL_0__11810_ (
);

FILL FILL227240x276640 (
);

AND2X2 _19432_ (
    .A(_8323_),
    .B(_8322_),
    .Y(_8320_[1])
);

AND2X2 _19012_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_7913_)
);

FILL FILL_0__9668_ (
);

OR2X2 _11939_ (
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .Y(_1849_)
);

AND2X2 _11519_ (
    .A(_1584_),
    .B(_1583_),
    .Y(_1521_[31])
);

FILL FILL_1_BUFX2_insert101 (
);

FILL FILL386080x98800 (
);

FILL FILL_1_BUFX2_insert103 (
);

FILL FILL_1_BUFX2_insert105 (
);

OR2X2 _15772_ (
    .A(_4720_),
    .B(_4721_),
    .Y(_4722_)
);

FILL FILL_0__15487_ (
);

FILL FILL_0__15067_ (
);

OR2X2 _15352_ (
    .A(_4308_),
    .B(_4293_),
    .Y(_4309_)
);

FILL FILL_1__8624_ (
);

FILL FILL468920x123500 (
);

FILL FILL414200x69160 (
);

FILL FILL_1__14807_ (
);

FILL FILL430920x44460 (
);

AND2X2 _16977_ (
    .A(_4195__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_5908_)
);

AND2X2 _16557_ (
    .A(_4223__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_5495_)
);

FILL FILL363280x172900 (
);

OR2X2 _16137_ (
    .A(_5080_),
    .B(_5073_),
    .Y(_5081_)
);

OR2X2 _11692_ (
    .A(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .B(_1718__bF$buf3),
    .Y(_1660_)
);

FILL FILL_1__18640_ (
);

DFFSR _11272_ (
    .CLK(clk_bF$buf5),
    .D(_1389_[10]),
    .Q(\datapath_1.regfile_1.regOut[22] [10]),
    .R(rst_bF$buf112),
    .S(vdd)
);

FILL FILL_0__17633_ (
);

FILL FILL_0__17213_ (
);

FILL FILL485640x360620 (
);

OR2X2 _8899_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .B(_266__bF$buf4),
    .Y(_238_)
);

FILL FILL293360x177840 (
);

OR2X2 _8479_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .B(_68__bF$buf2),
    .Y(_18_)
);

FILL FILL14440x14820 (
);

FILL FILL101840x167960 (
);

FILL FILL_1__10307_ (
);

FILL FILL219640x291460 (
);

OR2X2 _9840_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_725_)
);

OR2X2 _9420_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_505_)
);

OR2X2 _9000_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_285_)
);

NAND3X1 _12897_ (
    .A(_2279_),
    .B(\datapath_1.alu_1.ALUInA [18]),
    .C(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2462_)
);

FILL FILL_1__19425_ (
);

OR2X2 _12477_ (
    .A(_2056_),
    .B(_2069_),
    .Y(_2070_)
);

DFFSR _12057_ (
    .CLK(clk_bF$buf1),
    .D(_1785_[21]),
    .Q(\datapath_1.regfile_1.regOut[28] [21]),
    .R(rst_bF$buf62),
    .S(vdd)
);

FILL FILL_1__14140_ (
);

FILL FILL418000x69160 (
);

AND2X2 _18703_ (
    .A(_6232__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_7609_)
);

FILL FILL_0__13973_ (
);

FILL FILL342000x256880 (
);

FILL FILL_0__8939_ (
);

FILL FILL52440x306280 (
);

FILL FILL_1__15765_ (
);

FILL FILL_1__15345_ (
);

FILL FILL437760x281580 (
);

FILL FILL356440x217360 (
);

FILL FILL_1__10060_ (
);

FILL FILL_0__14758_ (
);

DFFSR _14623_ (
    .CLK(clk_bF$buf42),
    .D(_3738_[29]),
    .Q(\control_1.op [3]),
    .R(rst_bF$buf100),
    .S(vdd)
);

OR2X2 _14203_ (
    .A(MemToReg_bF$buf3),
    .B(ALUOut[20]),
    .Y(_3580_)
);

OR2X2 _17095_ (
    .A(_6023_),
    .B(_6022_),
    .Y(_6024_)
);

FILL FILL_0__18591_ (
);

FILL FILL274360x123500 (
);

FILL FILL_0__18171_ (
);

FILL FILL38000x29640 (
);

FILL FILL107920x158080 (
);

AND2X2 _15828_ (
    .A(_4187__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_4777_)
);

AND2X2 _15408_ (
    .A(_4217__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_4364_)
);

FILL FILL213560x232180 (
);

OR2X2 _10963_ (
    .A(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .B(_1322__bF$buf0),
    .Y(_1294_)
);

FILL FILL_0__10678_ (
);

OR2X2 _10543_ (
    .A(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .B(_1124__bF$buf4),
    .Y(_1074_)
);

DFFSR _10123_ (
    .CLK(clk_bF$buf74),
    .D(_795_[22]),
    .Q(\datapath_1.regfile_1.regOut[13] [22]),
    .R(rst_bF$buf105),
    .S(vdd)
);

FILL FILL_0__16904_ (
);

FILL FILL185440x286520 (
);

FILL FILL_0__19376_ (
);

AND2X2 _19241_ (
    .A(_6216__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_8138_)
);

FILL FILL_0__14091_ (
);

FILL FILL_0__9897_ (
);

FILL FILL272080x197600 (
);

FILL FILL_0__9057_ (
);

OR2X2 _11748_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_1697_)
);

OR2X2 _11328_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_1477_)
);

FILL FILL_0__12404_ (
);

FILL FILL117040x247000 (
);

FILL FILL_0__15296_ (
);

AND2X2 _15581_ (
    .A(_4195__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_4534_)
);

FILL FILL34200x281580 (
);

FILL FILL421040x182780 (
);

NOR3X1 _15161_ (
    .A(_4121_),
    .B(_4004_),
    .C(_4123_),
    .Y(\datapath_1.regfile_1.regEn [27])
);

FILL FILL_0__13609_ (
);

FILL FILL_1__17088_ (
);

AND2X2 _16786_ (
    .A(_4146__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_5720_)
);

OR2X2 _16366_ (
    .A(_5305_),
    .B(_5306_),
    .Y(_5307_)
);

FILL FILL79800x79040 (
);

FILL FILL96520x29640 (
);

AND2X2 _11081_ (
    .A(_1352_),
    .B(_1351_),
    .Y(_1323_[14])
);

FILL FILL_0__17862_ (
);

FILL FILL433200x39520 (
);

OR2X2 _12286_ (
    .A(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .B(_1982__bF$buf3),
    .Y(_1976_)
);

FILL FILL288040x326040 (
);

FILL FILL_0__18647_ (
);

OR2X2 _18932_ (
    .A(_7830_),
    .B(_7833_),
    .Y(_7834_)
);

FILL FILL_0__18227_ (
);

OR2X2 _18512_ (
    .A(_7405_),
    .B(_7420_),
    .Y(_7421_)
);

FILL FILL_0__13362_ (
);

FILL FILL_0__8748_ (
);

FILL FILL_1__9391_ (
);

FILL FILL_1__15994_ (
);

DFFSR _14852_ (
    .CLK(clk_bF$buf38),
    .D(_3870_[0]),
    .Q(_2_[0]),
    .R(rst_bF$buf15),
    .S(vdd)
);

FILL FILL_0__14567_ (
);

OR2X2 _14432_ (
    .A(vdd),
    .B(\datapath_1.Data [21]),
    .Y(_3714_)
);

AND2X2 _14012_ (
    .A(_3350__bF$buf0),
    .B(_2_[13]),
    .Y(_3430_)
);

FILL FILL109440x128440 (
);

AND2X2 _15637_ (
    .A(_4135__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_4589_)
);

AND2X2 _15217_ (
    .A(_4169_),
    .B(_4139_),
    .Y(_4175_)
);

FILL FILL471960x24700 (
);

DFFSR _10772_ (
    .CLK(clk_bF$buf109),
    .D(_1125_[26]),
    .Q(\datapath_1.regfile_1.regOut[18] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

FILL FILL_0__10067_ (
);

AND2X2 _10352_ (
    .A(_986_),
    .B(_985_),
    .Y(_927_[29])
);

FILL FILL_0__16713_ (
);

FILL FILL186200x0 (
);

FILL FILL264480x24700 (
);

FILL FILL87400x83980 (
);

OR2X2 _19470_ (
    .A(gnd),
    .B(_8385__bF$buf1),
    .Y(_8349_)
);

FILL FILL_0__19185_ (
);

OR2X2 _19050_ (
    .A(_7949_),
    .B(_7945_),
    .Y(_7950_)
);

FILL FILL66120x4940 (
);

OR2X2 _8920_ (
    .A(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .B(_266__bF$buf2),
    .Y(_252_)
);

OR2X2 _8500_ (
    .A(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .B(_68__bF$buf1),
    .Y(_32_)
);

FILL FILL_0__9286_ (
);

OR2X2 _11977_ (
    .A(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .B(_1850__bF$buf1),
    .Y(_1810_)
);

FILL FILL_1__18925_ (
);

OR2X2 _11557_ (
    .A(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .B(_1652__bF$buf2),
    .Y(_1590_)
);

FILL FILL_1__18505_ (
);

DFFSR _11137_ (
    .CLK(clk_bF$buf51),
    .D(_1323_[4]),
    .Q(\datapath_1.regfile_1.regOut[21] [4]),
    .R(rst_bF$buf12),
    .S(vdd)
);

FILL FILL353400x251940 (
);

FILL FILL27360x128440 (
);

FILL FILL_0__12633_ (
);

FILL FILL_0__12213_ (
);

AND2X2 _15390_ (
    .A(_4154__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_4346_)
);

OR2X2 _9705_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_655_)
);

FILL FILL_1__8662_ (
);

FILL FILL471200x148200 (
);

FILL FILL_1__14425_ (
);

FILL FILL_1__14005_ (
);

FILL FILL370120x167960 (
);

FILL FILL_0__13838_ (
);

AND2X2 _13703_ (
    .A(_3081__bF$buf2),
    .B(ALUOut[16]),
    .Y(_3182_)
);

FILL FILL454480x123500 (
);

FILL FILL495520x39520 (
);

OR2X2 _16595_ (
    .A(_5531_),
    .B(_5530_),
    .Y(_5532_)
);

OR2X2 _16175_ (
    .A(_5118_),
    .B(_5115_),
    .Y(_5119_)
);

FILL FILL278920x375440 (
);

FILL FILL93480x163020 (
);

FILL FILL101840x237120 (
);

FILL FILL288040x39520 (
);

FILL FILL_0__17251_ (
);

FILL FILL183920x335920 (
);

AND2X2 _14908_ (
    .A(_3951_),
    .B(_3950_),
    .Y(_3936_[7])
);

FILL FILL11400x123500 (
);

AND2X2 _12095_ (
    .A(_1868_),
    .B(_1867_),
    .Y(_1851_[8])
);

FILL FILL_0__18876_ (
);

FILL FILL392160x54340 (
);

AND2X2 _18741_ (
    .A(_6282__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[0] [21]),
    .Y(_7646_)
);

FILL FILL_0__18456_ (
);

AND2X2 _18321_ (
    .A(_6323__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_7232_)
);

FILL FILL_0__18036_ (
);

FILL FILL_0__13591_ (
);

FILL FILL482600x93860 (
);

FILL FILL_0__8977_ (
);

FILL FILL414200x365560 (
);

OR2X2 _10828_ (
    .A(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .B(_1256__bF$buf2),
    .Y(_1224_)
);

OR2X2 _10408_ (
    .A(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .B(_1058__bF$buf4),
    .Y(_1004_)
);

FILL FILL_1__12911_ (
);

FILL FILL_0__11904_ (
);

FILL FILL_1__15383_ (
);

FILL FILL463600x163020 (
);

DFFSR _19526_ (
    .CLK(clk_bF$buf100),
    .D(_8320_[3]),
    .Q(\datapath_1.regfile_1.regOut[0] [3]),
    .R(rst_bF$buf68),
    .S(vdd)
);

OR2X2 _19106_ (
    .A(_8004_),
    .B(_8003_),
    .Y(_8005_)
);

OR2X2 _14661_ (
    .A(\datapath_1.rd1 [11]),
    .B(_3869__bF$buf4),
    .Y(_3827_)
);

FILL FILL_0__14376_ (
);

OR2X2 _14241_ (
    .A(\datapath_1.ALUResult [0]),
    .B(_3671__bF$buf0),
    .Y(_3607_)
);

FILL FILL241680x330980 (
);

FILL FILL323760x148200 (
);

AND2X2 _15866_ (
    .A(_4814_),
    .B(_4065__bF$buf7),
    .Y(\datapath_1.rd2 [9])
);

OR2X2 _15446_ (
    .A(_4400_),
    .B(_4399_),
    .Y(_4401_)
);

AND2X2 _15026_ (
    .A(_4014_),
    .B(_4011_),
    .Y(_4015_)
);

OR2X2 _10581_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_1099_)
);

OR2X2 _10161_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_879_)
);

FILL FILL285000x360620 (
);

FILL FILL_0__16102_ (
);

FILL FILL399000x108680 (
);

FILL FILL266000x197600 (
);

DFFSR _11786_ (
    .CLK(clk_bF$buf84),
    .D(_1653_[8]),
    .Q(\datapath_1.regfile_1.regOut[26] [8]),
    .R(rst_bF$buf11),
    .S(vdd)
);

AND2X2 _11366_ (
    .A(_1502_),
    .B(_1501_),
    .Y(_1455_[23])
);

FILL FILL_0__17727_ (
);

FILL FILL_0__12862_ (
);

FILL FILL_0__12022_ (
);

FILL FILL76760x340860 (
);

OR2X2 _9934_ (
    .A(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .B(_794__bF$buf3),
    .Y(_768_)
);

OR2X2 _9514_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .B(_596__bF$buf2),
    .Y(_548_)
);

FILL FILL_1__8471_ (
);

FILL FILL116280x108680 (
);

FILL FILL_1__14234_ (
);

AND2X2 _13932_ (
    .A(_3344__bF$buf3),
    .B(vdd),
    .Y(_3361_)
);

FILL FILL_0__13227_ (
);

AND2X2 _13512_ (
    .A(_3029_),
    .B(_3028_),
    .Y(_1_[7])
);

FILL FILL254600x291460 (
);

FILL FILL234080x326040 (
);

FILL FILL_1__9676_ (
);

BUFX2 BUFX2_insert1060 (
    .A(_4241_),
    .Y(_4241__bF$buf4)
);

FILL FILL429400x330980 (
);

BUFX2 BUFX2_insert1061 (
    .A(_4241_),
    .Y(_4241__bF$buf3)
);

FILL FILL_0__17480_ (
);

BUFX2 BUFX2_insert1062 (
    .A(_4241_),
    .Y(_4241__bF$buf2)
);

BUFX2 BUFX2_insert1063 (
    .A(_4241_),
    .Y(_4241__bF$buf1)
);

BUFX2 BUFX2_insert1064 (
    .A(_4241_),
    .Y(_4241__bF$buf0)
);

BUFX2 BUFX2_insert1065 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf4 )
);

BUFX2 BUFX2_insert1066 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf3 )
);

FILL FILL_1__15859_ (
);

BUFX2 BUFX2_insert1067 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf2 )
);

BUFX2 BUFX2_insert1068 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf1 )
);

BUFX2 BUFX2_insert1069 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf0 )
);

FILL FILL_1__10994_ (
);

OR2X2 _14717_ (
    .A(vdd),
    .B(\datapath_1.a [30]),
    .Y(_3864_)
);

FILL FILL218120x34580 (
);

BUFX2 BUFX2_insert880 (
    .A(_398_),
    .Y(_398__bF$buf2)
);

BUFX2 BUFX2_insert881 (
    .A(_398_),
    .Y(_398__bF$buf1)
);

FILL FILL137560x360620 (
);

BUFX2 BUFX2_insert882 (
    .A(_398_),
    .Y(_398__bF$buf0)
);

BUFX2 BUFX2_insert883 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf4 )
);

BUFX2 BUFX2_insert884 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf3 )
);

BUFX2 BUFX2_insert885 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf2 )
);

BUFX2 BUFX2_insert886 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf1 )
);

AND2X2 _17189_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_6117_)
);

BUFX2 BUFX2_insert887 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf0 )
);

BUFX2 BUFX2_insert888 (
    .A(_3671_),
    .Y(_3671__bF$buf4)
);

BUFX2 BUFX2_insert889 (
    .A(_3671_),
    .Y(_3671__bF$buf3)
);

FILL FILL323760x375440 (
);

FILL FILL_0__18685_ (
);

AND2X2 _18970_ (
    .A(_7871_),
    .B(_4065__bF$buf1),
    .Y(\datapath_1.rd1 [24])
);

AND2X2 _18550_ (
    .A(_6255__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_7458_)
);

AND2X2 _18130_ (
    .A(_6206__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_7044_)
);

FILL FILL145160x19760 (
);

FILL FILL_0__8786_ (
);

DFFSR _10637_ (
    .CLK(clk_bF$buf27),
    .D(_1059_[20]),
    .Q(\datapath_1.regfile_1.regOut[17] [20]),
    .R(rst_bF$buf28),
    .S(vdd)
);

AND2X2 _10217_ (
    .A(_916_),
    .B(_915_),
    .Y(_861_[27])
);

FILL FILL463600x256880 (
);

FILL FILL_0__11713_ (
);

FILL FILL355680x350740 (
);

AND2X2 _19335_ (
    .A(_6312__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_8231_)
);

AND2X2 _14890_ (
    .A(_3939_),
    .B(_3938_),
    .Y(_3936_[1])
);

FILL FILL_0__14185_ (
);

DFFSR _14470_ (
    .CLK(clk_bF$buf31),
    .D(_3672_[5]),
    .Q(\datapath_1.Data [5]),
    .R(rst_bF$buf85),
    .S(vdd)
);

OR2X2 _14050_ (
    .A(_3462_),
    .B(_3459_),
    .Y(\datapath_1.alu_1.ALUInB [18])
);

FILL FILL356440x19760 (
);

FILL FILL_0__12918_ (
);

AND2X2 _15675_ (
    .A(_4181__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[0] [7]),
    .Y(_4626_)
);

NOR3X1 _15255_ (
    .A(_4132_),
    .B(\datapath_1.PCJump [19]),
    .C(_4153_),
    .Y(_4213_)
);

DFFSR _10390_ (
    .CLK(clk_bF$buf100),
    .D(_927_[31]),
    .Q(\datapath_1.regfile_1.regOut[15] [31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

FILL FILL220400x365560 (
);

FILL FILL_0__16751_ (
);

FILL FILL_0__16331_ (
);

FILL FILL253080x34580 (
);

FILL FILL186960x69160 (
);

OR2X2 _11595_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_1615_)
);

OR2X2 _11175_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_1395_)
);

FILL FILL_0__17956_ (
);

OR2X2 _17821_ (
    .A(_6736_),
    .B(_6739_),
    .Y(_6740_)
);

AND2X2 _17401_ (
    .A(_6326__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_6327_)
);

FILL FILL_0__17116_ (
);

FILL FILL_0__12251_ (
);

FILL FILL353400x0 (
);

DFFSR _9743_ (
    .CLK(clk_bF$buf0),
    .D(_597_[29]),
    .Q(\datapath_1.regfile_1.regOut[10] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

AND2X2 _9323_ (
    .A(_460_),
    .B(_459_),
    .Y(_399_[30])
);

AND2X2 _18606_ (
    .A(_6293__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_7513_)
);

FILL FILL_0__13876_ (
);

FILL FILL_0__13456_ (
);

AND2X2 _13741_ (
    .A(_3087__bF$buf4),
    .B(\datapath_1.ALUResult [21]),
    .Y(_3215_)
);

FILL FILL_0__13036_ (
);

OR2X2 _13321_ (
    .A(_2848_),
    .B(_2861_),
    .Y(_2862_)
);

FILL FILL_1__9065_ (
);

OR2X2 _14946_ (
    .A(\datapath_1.mux_pcsrc.dout [20]),
    .B(_4001__bF$buf0),
    .Y(_3977_)
);

OR2X2 _14526_ (
    .A(memoryOutData[9]),
    .B(_3803__bF$buf0),
    .Y(_3757_)
);

OR2X2 _14106_ (
    .A(_3510_),
    .B(_3507_),
    .Y(\datapath_1.alu_1.ALUInB [26])
);

FILL FILL_0__15602_ (
);

FILL FILL68400x187720 (
);

FILL FILL208240x182780 (
);

FILL FILL_0__18074_ (
);

FILL FILL3040x4940 (
);

FILL FILL318440x49400 (
);

FILL FILL268280x296400 (
);

FILL FILL505400x316160 (
);

FILL FILL_1__11168_ (
);

FILL FILL_0__8595_ (
);

OR2X2 _10866_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_1249_)
);

OR2X2 _10446_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_1029_)
);

OR2X2 _10026_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_809_)
);

FILL FILL_0__11942_ (
);

FILL FILL_0__11102_ (
);

OR2X2 _19144_ (
    .A(_8039_),
    .B(_8042_),
    .Y(_8043_)
);

FILL FILL192280x9880 (
);

FILL FILL148200x370500 (
);

FILL FILL_1__13734_ (
);

FILL FILL158080x316160 (
);

FILL FILL_0__12727_ (
);

AND2X2 _15484_ (
    .A(_4210__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_4438_)
);

AND2X2 _15064_ (
    .A(_4052_),
    .B(_4041_),
    .Y(_4053_)
);

FILL FILL_1__8756_ (
);

FILL FILL175560x326040 (
);

FILL FILL_0__16980_ (
);

FILL FILL89680x54340 (
);

FILL FILL_1__14519_ (
);

FILL FILL161880x350740 (
);

FILL FILL155040x4940 (
);

FILL FILL271320x69160 (
);

AND2X2 _16689_ (
    .A(_4239__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_5625_)
);

AND2X2 _16269_ (
    .A(_4214__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_5211_)
);

FILL FILL9880x158080 (
);

FILL FILL256880x256880 (
);

FILL FILL_0__17765_ (
);

AND2X2 _17630_ (
    .A(_6247__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_6552_)
);

FILL FILL_0__17345_ (
);

AND2X2 _17210_ (
    .A(_6137_),
    .B(_4065__bF$buf4),
    .Y(\datapath_1.rd2 [30])
);

FILL FILL66120x370500 (
);

FILL FILL357200x335920 (
);

FILL FILL_0__12480_ (
);

FILL FILL446120x79040 (
);

FILL FILL169480x49400 (
);

FILL FILL_1__10439_ (
);

DFFSR _9972_ (
    .CLK(clk_bF$buf99),
    .D(_729_[0]),
    .Q(\datapath_1.regfile_1.regOut[12] [0]),
    .R(rst_bF$buf72),
    .S(vdd)
);

OR2X2 _9552_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_573_)
);

OR2X2 _9132_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_353_)
);

FILL FILL_1__19557_ (
);

DFFSR _12189_ (
    .CLK(clk_bF$buf105),
    .D(_1851_[24]),
    .Q(\datapath_1.regfile_1.regOut[29] [24]),
    .R(rst_bF$buf34),
    .S(vdd)
);

FILL FILL93480x326040 (
);

OR2X2 _18835_ (
    .A(_7735_),
    .B(_7738_),
    .Y(_7739_)
);

FILL FILL_0_BUFX2_insert521 (
);

AND2X2 _18415_ (
    .A(_6282__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_7325_)
);

FILL FILL_0_BUFX2_insert523 (
);

AND2X2 _13970_ (
    .A(_3350__bF$buf3),
    .B(_2_[7]),
    .Y(_3394_)
);

FILL FILL_0_BUFX2_insert524 (
);

FILL FILL_0__13685_ (
);

FILL FILL_0_BUFX2_insert525 (
);

OR2X2 _13550_ (
    .A(ALUOut[20]),
    .B(_3079__bF$buf2),
    .Y(_3055_)
);

AOI21X1 _13130_ (
    .A(_2547_),
    .B(_2682_),
    .C(_2675_),
    .Y(_2683_)
);

FILL FILL_0_BUFX2_insert526 (
);

FILL FILL_0_BUFX2_insert527 (
);

FILL FILL_0_BUFX2_insert529 (
);

FILL FILL397480x237120 (
);

FILL FILL54720x143260 (
);

FILL FILL_1__10192_ (
);

OR2X2 _14755_ (
    .A(_2_[0]),
    .B(vdd),
    .Y(_3934_)
);

AND2X2 _14335_ (
    .A(_3669_),
    .B(_3668_),
    .Y(_3606_[31])
);

FILL FILL446120x316160 (
);

FILL FILL_0__15831_ (
);

FILL FILL290320x306280 (
);

FILL FILL432440x340860 (
);

FILL FILL447640x88920 (
);

FILL FILL349600x350740 (
);

FILL FILL_1__17623_ (
);

OR2X2 _10675_ (
    .A(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .B(_1190__bF$buf3),
    .Y(_1142_)
);

DFFSR _10255_ (
    .CLK(clk_bF$buf93),
    .D(_861_[25]),
    .Q(\datapath_1.regfile_1.regOut[14] [25]),
    .R(rst_bF$buf41),
    .S(vdd)
);

FILL FILL_0__16616_ (
);

AND2X2 _16901_ (
    .A(_4200__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_5833_)
);

FILL FILL_0__11331_ (
);

FILL FILL430920x187720 (
);

OR2X2 _19373_ (
    .A(_8266_),
    .B(_8267_),
    .Y(_8268_)
);

FILL FILL_0__19088_ (
);

DFFSR _8823_ (
    .CLK(clk_bF$buf102),
    .D(_135_[12]),
    .Q(\datapath_1.regfile_1.regOut[3] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

BUFX2 _8403_ (
    .A(_1_[11]),
    .Y(memoryAddress[11])
);

FILL FILL115520x163020 (
);

FILL FILL408880x296400 (
);

FILL FILL_0__9189_ (
);

FILL FILL_1__13123_ (
);

FILL FILL180120x345800 (
);

FILL FILL_0__12956_ (
);

INVX1 _12821_ (
    .A(_2378_),
    .Y(_2386_)
);

FILL FILL_0__12536_ (
);

AND2X2 _12401_ (
    .A(_2032_),
    .B(_2031_),
    .Y(_1983_[24])
);

OR2X2 _15293_ (
    .A(_4248_),
    .B(_4249_),
    .Y(_4250_)
);

FILL FILL85880x207480 (
);

DFFSR _9608_ (
    .CLK(clk_bF$buf83),
    .D(_531_[23]),
    .Q(\datapath_1.regfile_1.regOut[9] [23]),
    .R(rst_bF$buf17),
    .S(vdd)
);

FILL FILL188480x365560 (
);

FILL FILL221160x103740 (
);

FILL FILL307040x118560 (
);

AND2X2 _13606_ (
    .A(_3084__bF$buf0),
    .B(\aluControl_1.inst [0]),
    .Y(_3099_)
);

OR2X2 _16498_ (
    .A(_5435_),
    .B(_5436_),
    .Y(_5437_)
);

AND2X2 _16078_ (
    .A(_4130__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_5023_)
);

FILL FILL_0__17994_ (
);

FILL FILL_0__17574_ (
);

FILL FILL_0__17154_ (
);

OR2X2 _9781_ (
    .A(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .B(_728__bF$buf4),
    .Y(_686_)
);

OR2X2 _9361_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(_530__bF$buf4),
    .Y(_466_)
);

FILL FILL_1__19366_ (
);

FILL FILL_0__10602_ (
);

FILL FILL356440x103740 (
);

OR2X2 _18644_ (
    .A(_7517_),
    .B(_7550_),
    .Y(_7551_)
);

AND2X2 _18224_ (
    .A(_6255__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_7137_)
);

FILL FILL319960x247000 (
);

FILL FILL_0__13494_ (
);

FILL FILL_0__13074_ (
);

FILL FILL119320x59280 (
);

FILL FILL195320x9880 (
);

FILL FILL_0__9401_ (
);

AND2X2 _19429_ (
    .A(_8321_),
    .B(_8384_),
    .Y(_8320_[0])
);

AND2X2 _19009_ (
    .A(_6297__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_7910_)
);

DFFSR _14984_ (
    .CLK(clk_bF$buf77),
    .D(_3936_[3]),
    .Q(\datapath_1.mux_iord.din0 [3]),
    .R(rst_bF$buf65),
    .S(vdd)
);

FILL FILL_0__14699_ (
);

FILL FILL_0__14279_ (
);

OR2X2 _14564_ (
    .A(IRWrite_bF$buf4),
    .B(\datapath_1.PCJump [24]),
    .Y(_3782_)
);

OR2X2 _14144_ (
    .A(\datapath_1.Data [0]),
    .B(_3605__bF$buf2),
    .Y(_3541_)
);

FILL FILL6840x192660 (
);

FILL FILL_0__15220_ (
);

OR2X2 _15769_ (
    .A(_4703_),
    .B(_4718_),
    .Y(_4719_)
);

OR2X2 _15349_ (
    .A(_4304_),
    .B(_4305_),
    .Y(_4306_)
);

FILL FILL130720x222300 (
);

AND2X2 _10484_ (
    .A(_1054_),
    .B(_1053_),
    .Y(_993_[30])
);

AND2X2 _10064_ (
    .A(_834_),
    .B(_833_),
    .Y(_795_[19])
);

FILL FILL_1__17012_ (
);

FILL FILL_0__16845_ (
);

FILL FILL_0__16425_ (
);

AND2X2 _16710_ (
    .A(_4154__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_5645_)
);

FILL FILL_0__11980_ (
);

FILL FILL_0__11560_ (
);

FILL FILL115520x256880 (
);

AND2X2 _19182_ (
    .A(_6247__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_8080_)
);

OR2X2 _8632_ (
    .A(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .B(_134__bF$buf2),
    .Y(_100_)
);

endmodule
